VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

VIA via1_2_560_340_1_1_300_300
  VIARULE Via1Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal1 via1 metal2 ;
  CUTSPACING 0.08 0.08 ;
  ENCLOSURE 0.105 0.05 0.035 0.035 ;
END via1_2_560_340_1_1_300_300

VIA via2_3_560_340_1_1_320_320
  VIARULE Via2Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal2 via2 metal3 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.035 0.035 ;
END via2_3_560_340_1_1_320_320

VIA via3_4_560_340_1_1_320_320
  VIARULE Via3Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal3 via3 metal4 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.035 0.035 ;
END via3_4_560_340_1_1_320_320

VIA via4_5_560_340_1_1_600_600
  VIARULE Via4Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal4 via4 metal5 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0 0 ;
END via4_5_560_340_1_1_600_600

VIA via5_6_560_340_1_1_600_600
  VIARULE Via5Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal5 via5 metal6 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0.07 0 ;
END via5_6_560_340_1_1_600_600

VIA via1_2_2400_340_1_8_300_300
  VIARULE Via1Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal1 via1 metal2 ;
  CUTSPACING 0.08 0.08 ;
  ENCLOSURE 0.04 0.05 0.035 0.035 ;
  ROWCOL 1 8 ;
END via1_2_2400_340_1_8_300_300

VIA via2_3_2400_920_3_7_320_320
  VIARULE Via2Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal2 via2 metal3 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.035 0.035 ;
  ROWCOL 3 7 ;
END via2_3_2400_920_3_7_320_320

VIA via3_4_2400_920_3_7_320_320
  VIARULE Via3Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal3 via3 metal4 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.035 0.035 ;
  ROWCOL 3 7 ;
END via3_4_2400_920_3_7_320_320

VIA via4_5_2400_920_2_4_600_600
  VIARULE Via4Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal4 via4 metal5 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0 0 ;
  ROWCOL 2 4 ;
END via4_5_2400_920_2_4_600_600

VIA via5_6_2400_1120_2_4_600_600
  VIARULE Via5Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal5 via5 metal6 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0 0 ;
  ROWCOL 2 4 ;
END via5_6_2400_1120_2_4_600_600

VIA via6_7_2400_1120_1_3_600_600
  VIARULE Via6Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal6 via6 metal7 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0.13 0.13 ;
  ROWCOL 1 3 ;
END via6_7_2400_1120_1_3_600_600

VIA via7_8_2400_1320_1_1_1680_1680
  VIARULE Via7Array-0 ;
  CUTSIZE 0.4 0.4 ;
  LAYERS metal7 via7 metal8 ;
  CUTSPACING 0.44 0.44 ;
  ENCLOSURE 0 0 0.4 0 ;
END via7_8_2400_1320_1_1_1680_1680

VIA via6_7_560_2400_3_1_600_600
  VIARULE Via6Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal6 via6 metal7 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0.07 0 0.13 0.23 ;
  ROWCOL 3 1 ;
END via6_7_560_2400_3_1_600_600

VIA via7_8_2400_2400_1_1_1680_1680
  VIARULE Via7Array-0 ;
  CUTSIZE 0.4 0.4 ;
  LAYERS metal7 via7 metal8 ;
  CUTSPACING 0.44 0.44 ;
  ENCLOSURE 0 0.4 0.4 0 ;
END via7_8_2400_2400_1_1_1680_1680

VIA via6_7_1120_2400_3_1_600_600
  VIARULE Via6Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal6 via6 metal7 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0.21 0.23 0.21 0.23 ;
  ROWCOL 3 1 ;
END via6_7_1120_2400_3_1_600_600

MACRO top
  FOREIGN top 0 0 ;
  CLASS BLOCK ;
  SIZE 200 BY 105 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  199.93 41.755 200 41.825 ;
    END
  END clk
  PIN din
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  29.7 104.93 29.77 105 ;
    END
  END din
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  199.93 72.835 200 72.905 ;
    END
  END enable
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  169.92 0 169.99 0.07 ;
    END
  END rst
  PIN spike
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  114.44 104.93 114.51 105 ;
    END
  END spike
  PIN x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  0.82 0 0.89 0.07 ;
    END
  END x[0]
  PIN x[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  127.74 0 127.81 0.07 ;
    END
  END x[10]
  PIN x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  43 0 43.07 0.07 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  156.62 104.93 156.69 105 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.955 0.07 32.025 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 63.035 0.07 63.105 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  198.8 104.93 198.87 105 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  85.18 0 85.25 0.07 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 94.395 0.07 94.465 ;
    END
  END x[7]
  PIN x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  71.88 104.93 71.95 105 ;
    END
  END x[8]
  PIN x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  199.93 10.395 200 10.465 ;
    END
  END x[9]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal7 ;
        RECT  0 90.8 200 92 ;
        RECT  0 70.8 200 72 ;
        RECT  0 50.8 200 52 ;
        RECT  0 30.8 200 32 ;
        RECT  0 10.8 200 12 ;
      LAYER metal8 ;
        RECT  189.97 0 191.17 105 ;
        RECT  169.97 0 171.17 105 ;
        RECT  149.97 0 151.17 105 ;
        RECT  129.97 0 131.17 105 ;
        RECT  109.97 0 111.17 105 ;
        RECT  89.97 0 91.17 105 ;
        RECT  69.97 0 71.17 105 ;
        RECT  49.97 0 51.17 105 ;
        RECT  29.97 0 31.17 105 ;
        RECT  9.97 0 11.17 105 ;
      LAYER metal6 ;
        RECT  195.43 0 195.71 105 ;
        RECT  95.43 0 95.71 105 ;
        RECT  4.43 0 4.71 105 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal7 ;
        RECT  0 100.8 200 102 ;
        RECT  0 80.8 200 82 ;
        RECT  0 60.8 200 62 ;
        RECT  0 40.8 200 42 ;
        RECT  0 20.8 200 22 ;
      LAYER metal8 ;
        RECT  179.97 0 181.17 105 ;
        RECT  159.97 0 161.17 105 ;
        RECT  139.97 0 141.17 105 ;
        RECT  119.97 0 121.17 105 ;
        RECT  99.97 0 101.17 105 ;
        RECT  79.97 0 81.17 105 ;
        RECT  59.97 0 61.17 105 ;
        RECT  39.97 0 41.17 105 ;
        RECT  19.97 0 21.17 105 ;
      LAYER metal6 ;
        RECT  195.99 0 196.27 105 ;
        RECT  95.99 0 96.27 105 ;
        RECT  4.99 0 5.27 105 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
     RECT  0.57 1.315 7.79 103.685 ;
     RECT  7.79 1.315 11.84 89.265 ;
     RECT  7.79 92.315 11.84 103.685 ;
     RECT  11.84 1.315 47.63 103.685 ;
     RECT  47.63 1.315 50.98 89.425 ;
     RECT  47.63 92.315 50.98 103.685 ;
     RECT  50.98 1.315 96.39 103.685 ;
     RECT  96.39 1.315 114.51 104.965 ;
     RECT  114.51 1.315 184.43 103.685 ;
     RECT  184.43 1.315 191.9 7.085 ;
     RECT  184.43 10.395 191.9 103.685 ;
     RECT  191.9 1.315 199.5 103.685 ;
     RECT  199.5 10.395 199.82 10.465 ;
     RECT  199.5 95.935 199.82 96.005 ;
    LAYER metal2 ;
     RECT  169.16 0 169.8 0.035 ;
     RECT  85.18 0.035 85.25 0.245 ;
     RECT  127.74 0.035 127.81 0.245 ;
     RECT  43 0.035 43.07 0.385 ;
     RECT  9.56 0.035 9.63 1.17 ;
     RECT  169.16 0.035 169.99 1.17 ;
     RECT  0.82 0.035 0.89 1.33 ;
     RECT  0.82 1.33 4.64 2.73 ;
     RECT  95.5 1.33 95.64 2.73 ;
     RECT  99.975 2.57 101.165 2.73 ;
     RECT  195.5 1.33 195.64 2.73 ;
     RECT  119.975 2.57 121.165 5.83 ;
     RECT  139.975 2.57 141.165 5.83 ;
     RECT  159.975 2.57 161.165 5.83 ;
     RECT  179.975 2.57 181.165 5.83 ;
     RECT  95.5 2.73 101.165 6.335 ;
     RECT  189.975 1.17 191.165 6.335 ;
     RECT  143.32 6.335 144.91 6.405 ;
     RECT  109.975 1.17 111.165 7.23 ;
     RECT  169.16 1.17 171.165 7.23 ;
     RECT  189.49 6.335 191.165 7.23 ;
     RECT  19.975 2.57 21.165 8.63 ;
     RECT  39.975 2.57 41.165 8.63 ;
     RECT  59.975 2.57 61.165 8.63 ;
     RECT  79.975 2.57 81.165 8.63 ;
     RECT  95.5 6.335 101.59 9.135 ;
     RECT  95.5 9.135 102.54 9.94 ;
     RECT  149.975 1.17 151.165 9.94 ;
     RECT  169.16 7.23 169.99 9.94 ;
     RECT  184.36 8.995 184.43 9.94 ;
     RECT  49.975 1.17 51.165 9.975 ;
     RECT  9.56 1.17 11.165 10.03 ;
     RECT  29.975 1.17 31.165 10.03 ;
     RECT  49.975 9.975 53.9 10.03 ;
     RECT  69.975 1.17 71.165 10.03 ;
     RECT  89.975 1.17 91.165 10.03 ;
     RECT  53.83 10.03 53.9 10.395 ;
     RECT  195.5 2.73 196.2 10.395 ;
     RECT  53.83 10.395 57.13 10.465 ;
     RECT  9.56 10.03 9.82 10.535 ;
     RECT  129.975 1.17 131.165 10.815 ;
     RECT  144.84 6.405 144.91 10.815 ;
     RECT  149.975 9.94 152.89 10.815 ;
     RECT  119.95 9.94 121.54 10.955 ;
     RECT  129.64 10.815 132.94 10.955 ;
     RECT  136.86 9.135 136.93 10.955 ;
     RECT  144.84 10.815 152.89 10.955 ;
     RECT  162.13 10.815 162.2 10.955 ;
     RECT  95.5 9.94 105.77 11.095 ;
     RECT  119.76 10.955 121.54 11.095 ;
     RECT  160.04 10.955 162.2 11.095 ;
     RECT  189.49 7.23 189.56 11.095 ;
     RECT  95.5 11.095 107.29 11.27 ;
     RECT  126.41 10.955 136.93 11.27 ;
     RECT  168.02 9.94 169.99 11.27 ;
     RECT  183.6 9.94 184.43 11.27 ;
     RECT  144.84 10.955 155.36 11.515 ;
     RECT  159.85 11.095 162.58 11.515 ;
     RECT  116.91 11.095 121.54 11.655 ;
     RECT  126.41 11.27 140.68 11.655 ;
     RECT  144.84 11.515 162.58 11.655 ;
     RECT  168.02 11.27 170.68 11.655 ;
     RECT  180.22 11.27 184.43 11.655 ;
     RECT  95.5 11.27 110.68 11.725 ;
     RECT  116.91 11.655 162.58 11.795 ;
     RECT  167.07 11.655 170.68 11.795 ;
     RECT  53.83 10.465 55.8 11.865 ;
     RECT  115.01 11.795 170.68 11.935 ;
     RECT  180.22 11.655 184.62 11.935 ;
     RECT  189.49 11.095 189.94 11.935 ;
     RECT  115.01 11.935 172.08 12.215 ;
     RECT  107.22 11.725 110.68 12.355 ;
     RECT  114.82 12.215 172.08 12.355 ;
     RECT  107.22 12.355 172.08 12.67 ;
     RECT  177.9 11.935 189.94 12.67 ;
     RECT  9.75 10.535 9.82 14.735 ;
     RECT  95.5 11.725 102.54 14.735 ;
     RECT  9.56 14.735 9.82 14.98 ;
     RECT  39.58 9.135 39.65 14.98 ;
     RECT  39.58 14.98 41.17 15.015 ;
     RECT  68.46 14.98 68.72 15.015 ;
     RECT  39.58 15.015 42.69 15.155 ;
     RECT  87.08 11.795 87.15 15.17 ;
     RECT  94.68 14.735 102.54 15.17 ;
     RECT  39.58 15.155 44.78 15.855 ;
     RECT  67.89 15.015 68.72 15.855 ;
     RECT  66.75 15.855 72.33 15.995 ;
     RECT  25.14 10.395 25.21 16.135 ;
     RECT  31.03 15.855 34.71 16.135 ;
     RECT  66.56 15.995 72.33 16.135 ;
     RECT  23.62 16.135 34.71 16.31 ;
     RECT  53.83 11.865 54.09 16.31 ;
     RECT  60.86 16.135 72.33 16.31 ;
     RECT  15.22 16.31 15.68 16.695 ;
     RECT  39.58 15.855 48.2 16.695 ;
     RECT  60.86 16.31 75.68 16.695 ;
     RECT  82.14 14.98 82.97 16.695 ;
     RECT  9.56 14.98 11.15 16.765 ;
     RECT  15.22 16.695 19.13 16.835 ;
     RECT  23.62 16.31 35.68 16.835 ;
     RECT  39.58 16.695 49.72 16.835 ;
     RECT  53.83 16.31 55.68 16.835 ;
     RECT  15.22 16.835 35.68 16.975 ;
     RECT  39.58 16.835 55.68 16.975 ;
     RECT  60.86 16.695 82.97 16.975 ;
     RECT  15.22 16.975 82.97 17.535 ;
     RECT  87.08 15.17 102.54 18.43 ;
     RECT  15.22 17.535 83.16 18.585 ;
     RECT  107.22 12.67 189.94 18.655 ;
     RECT  94.68 18.43 102.54 19.075 ;
     RECT  106.46 18.655 189.94 19.075 ;
     RECT  15.22 18.585 82.59 21.595 ;
     RECT  14.69 21.595 82.59 22.575 ;
     RECT  87.08 18.43 87.15 22.575 ;
     RECT  14.69 22.575 87.15 22.715 ;
     RECT  14.12 22.715 87.15 23.57 ;
     RECT  94.68 19.075 189.94 23.57 ;
     RECT  9.56 16.765 9.82 23.695 ;
     RECT  14.12 23.57 189.94 23.695 ;
     RECT  9.56 23.695 189.94 29.645 ;
     RECT  9.56 29.645 188.99 29.785 ;
     RECT  106.46 29.785 188.99 29.925 ;
     RECT  106.65 29.925 188.99 31.605 ;
     RECT  0.82 2.73 5.2 31.955 ;
     RECT  9.56 29.785 102.54 32.865 ;
     RECT  89.975 32.865 102.54 33.775 ;
     RECT  106.65 31.605 188.23 33.775 ;
     RECT  89.975 33.775 188.23 35.525 ;
     RECT  106.84 35.525 188.23 35.875 ;
     RECT  106.84 35.875 189.18 36.855 ;
     RECT  9.56 32.865 84.87 36.925 ;
     RECT  89.975 35.525 102.54 38.03 ;
     RECT  10.7 36.925 84.87 39.165 ;
     RECT  94.11 38.03 102.54 40.355 ;
     RECT  106.84 36.855 189.37 40.355 ;
     RECT  195.5 10.395 199.82 41.825 ;
     RECT  94.11 40.355 189.37 43.17 ;
     RECT  89.975 43.17 189.37 43.575 ;
     RECT  10.89 39.165 84.87 47.355 ;
     RECT  10.7 47.355 84.87 48.195 ;
     RECT  89.975 43.575 188.99 49.23 ;
     RECT  90.69 49.23 188.99 52.675 ;
     RECT  90.69 52.675 189.18 54.37 ;
     RECT  89.975 54.37 189.18 57.63 ;
     RECT  90.69 57.63 189.18 58.205 ;
     RECT  91.45 58.205 189.18 58.275 ;
     RECT  9.75 48.195 84.87 61.985 ;
     RECT  91.45 58.275 188.99 62.77 ;
     RECT  89.975 62.77 188.99 63.875 ;
     RECT  9.75 61.985 83.73 66.675 ;
     RECT  89.975 63.875 189.56 66.675 ;
     RECT  9.75 66.675 189.56 67.935 ;
     RECT  9.75 67.935 189.75 68.005 ;
     RECT  9.75 68.005 91.165 68.83 ;
     RECT  195.5 41.825 196.2 72.835 ;
     RECT  9.75 68.83 87.34 73.97 ;
     RECT  9.75 73.97 91.165 75.845 ;
     RECT  14.12 75.845 91.165 75.985 ;
     RECT  15.22 75.985 91.165 80.03 ;
     RECT  15.22 80.03 87.34 81.095 ;
     RECT  9.75 75.845 9.82 82.915 ;
     RECT  14.69 81.095 87.34 82.915 ;
     RECT  95.5 68.005 189.75 83.125 ;
     RECT  95.5 83.125 188.99 83.545 ;
     RECT  9.75 82.915 87.34 83.825 ;
     RECT  9.75 83.825 9.82 83.965 ;
     RECT  9.56 83.965 9.82 84.035 ;
     RECT  14.31 83.825 87.34 84.525 ;
     RECT  15.22 84.525 87.34 85.17 ;
     RECT  95.5 83.545 188.61 87.535 ;
     RECT  95.5 87.535 188.99 87.605 ;
     RECT  15.22 85.17 91.165 88.375 ;
     RECT  14.88 88.375 91.165 88.43 ;
     RECT  0.06 31.955 5.2 88.445 ;
     RECT  95.5 87.605 189.18 88.935 ;
     RECT  14.88 88.43 87.34 89.25 ;
     RECT  14.88 89.25 41.55 89.425 ;
     RECT  46.04 89.25 87.34 89.425 ;
     RECT  14.88 89.425 16.85 89.565 ;
     RECT  21.34 89.425 28.82 89.565 ;
     RECT  46.04 89.425 55.23 89.565 ;
     RECT  79.86 89.425 87.34 89.565 ;
     RECT  9.56 84.035 9.63 89.635 ;
     RECT  14.88 89.565 14.95 89.635 ;
     RECT  22.48 89.565 26.54 89.705 ;
     RECT  35.97 89.425 41.55 89.705 ;
     RECT  53.07 89.565 55.23 89.705 ;
     RECT  26.09 89.705 26.54 89.845 ;
     RECT  46.99 89.565 47.06 89.845 ;
     RECT  53.26 89.705 55.23 89.845 ;
     RECT  60.29 89.425 75.56 89.845 ;
     RECT  81.57 89.565 87.34 89.845 ;
     RECT  26.28 89.845 26.54 89.98 ;
     RECT  39.77 89.705 41.55 89.98 ;
     RECT  9.56 89.635 14.95 89.985 ;
     RECT  26.47 89.98 26.54 89.985 ;
     RECT  40.72 89.98 41.55 90.125 ;
     RECT  75.49 89.845 75.56 90.265 ;
     RECT  69.6 89.845 71.165 90.405 ;
     RECT  0.06 88.445 0.13 90.545 ;
     RECT  84.04 89.845 87.34 90.545 ;
     RECT  95.5 88.935 189.37 91.945 ;
     RECT  95.5 91.945 110.68 92.085 ;
     RECT  110.22 92.085 110.68 92.61 ;
     RECT  115.01 91.945 189.37 92.61 ;
     RECT  115.01 92.61 128.95 93.205 ;
     RECT  133.82 92.61 189.37 93.205 ;
     RECT  141.99 93.205 175.88 93.485 ;
     RECT  87.08 90.545 87.34 93.57 ;
     RECT  115.22 93.205 128.95 94.01 ;
     RECT  185.22 93.205 189.37 94.01 ;
     RECT  115.77 94.01 128.95 94.185 ;
     RECT  173.91 93.485 175.88 94.185 ;
     RECT  126.22 94.185 127.43 94.325 ;
     RECT  133.82 93.205 137.5 94.325 ;
     RECT  141.99 93.485 168.85 94.325 ;
     RECT  179.8 93.205 181.39 94.325 ;
     RECT  117.48 94.185 122.11 94.465 ;
     RECT  127.36 94.325 127.43 94.465 ;
     RECT  149.21 94.325 154.6 94.465 ;
     RECT  158.9 94.325 168.28 94.465 ;
     RECT  173.91 94.185 173.98 94.465 ;
     RECT  55.16 89.845 55.23 94.605 ;
     RECT  141.99 94.325 144.91 94.605 ;
     RECT  149.21 94.465 154.03 94.605 ;
     RECT  95.5 92.085 102.92 94.745 ;
     RECT  159.975 94.465 168.28 94.885 ;
     RECT  117.48 94.465 121.165 94.94 ;
     RECT  149.21 94.605 149.85 94.94 ;
     RECT  179.975 94.325 181.39 94.94 ;
     RECT  41.48 90.125 41.55 94.97 ;
     RECT  159.975 94.885 165.43 95.165 ;
     RECT  39.975 94.97 41.55 95.865 ;
     RECT  118.24 94.94 121.165 95.865 ;
     RECT  133.82 94.325 133.89 95.865 ;
     RECT  189.3 94.01 189.37 96.005 ;
     RECT  195.5 72.835 199.82 96.005 ;
     RECT  19.975 94.97 21.165 98.23 ;
     RECT  39.975 95.865 41.165 98.23 ;
     RECT  59.975 94.97 61.165 98.23 ;
     RECT  79.975 94.97 81.165 98.23 ;
     RECT  95.5 94.745 101.59 98.23 ;
     RECT  119.975 95.865 121.165 98.23 ;
     RECT  139.975 97.77 141.165 98.23 ;
     RECT  159.975 95.165 161.165 98.23 ;
     RECT  179.975 94.94 181.165 98.23 ;
     RECT  101.52 98.23 101.59 98.805 ;
     RECT  146.93 98.735 147.38 98.805 ;
     RECT  9.56 89.985 11.165 99.63 ;
     RECT  29.975 93.57 31.165 99.63 ;
     RECT  49.975 93.57 51.165 99.63 ;
     RECT  69.975 90.405 71.165 99.63 ;
     RECT  87.08 93.57 91.165 99.63 ;
     RECT  109.975 99.17 111.165 99.63 ;
     RECT  129.975 99.17 131.165 99.63 ;
     RECT  149.975 99.17 151.165 99.63 ;
     RECT  169.975 99.17 171.165 99.63 ;
     RECT  189.975 99.17 191.165 99.63 ;
     RECT  4.5 88.445 5.2 102.27 ;
     RECT  95.5 98.23 96.46 102.27 ;
     RECT  195.5 96.005 196.2 102.27 ;
     RECT  47.75 102.795 48.77 102.865 ;
     RECT  48.32 102.865 48.77 103.005 ;
     RECT  87.08 99.63 87.15 103.005 ;
     RECT  96.06 102.27 96.46 103.37 ;
     RECT  5.06 102.27 5.2 103.67 ;
     RECT  96.06 103.37 101.165 103.67 ;
     RECT  196.06 102.27 196.2 103.67 ;
     RECT  19.975 103.37 21.165 103.83 ;
     RECT  39.975 103.37 41.165 103.83 ;
     RECT  59.975 103.37 61.165 103.83 ;
     RECT  79.975 103.37 81.165 103.83 ;
     RECT  96.39 103.67 101.165 103.83 ;
     RECT  119.975 103.37 121.165 103.83 ;
     RECT  139.975 103.37 141.165 103.83 ;
     RECT  159.975 103.37 161.165 103.83 ;
     RECT  179.975 103.37 181.165 103.83 ;
     RECT  9.56 99.63 9.63 104.965 ;
     RECT  29.7 102.795 29.77 104.965 ;
     RECT  71.88 104.755 71.95 104.965 ;
     RECT  96.39 103.83 96.46 104.965 ;
     RECT  114.44 104.755 114.51 104.965 ;
     RECT  156.62 104.755 156.69 104.965 ;
     RECT  198.8 104.755 198.87 104.965 ;
    LAYER metal3 ;
     RECT  0.035 31.955 0.13 32.025 ;
     RECT  0.035 94.395 0.13 94.465 ;
     RECT  0.035 63.035 0.69 63.105 ;
     RECT  0.06 90.475 0.82 90.545 ;
     RECT  0.82 88.375 4.5 90.545 ;
     RECT  4.5 1.33 4.64 102.27 ;
     RECT  4.64 2.73 5.06 102.27 ;
     RECT  5.06 2.73 5.2 103.67 ;
     RECT  9.75 25.515 9.88 25.585 ;
     RECT  9.56 36.855 9.88 36.925 ;
     RECT  9.75 48.195 9.88 48.265 ;
     RECT  9.58 58.135 9.88 58.205 ;
     RECT  9.86 68.915 9.88 68.985 ;
     RECT  9.88 25.515 9.95 26.985 ;
     RECT  9.95 26.215 10.01 26.985 ;
     RECT  9.56 0.035 10.02 0.105 ;
     RECT  9.88 79.135 10.21 79.765 ;
     RECT  9.88 58.135 10.89 58.625 ;
     RECT  10.89 53.235 11.08 53.305 ;
     RECT  10.89 58.135 11.08 60.305 ;
     RECT  10.02 0.035 11.12 10.03 ;
     RECT  10.02 93.57 11.12 99.63 ;
     RECT  11.08 57.855 11.27 60.445 ;
     RECT  11.27 33.635 11.46 33.705 ;
     RECT  9.88 36.855 11.46 37.625 ;
     RECT  11.27 42.455 11.46 42.525 ;
     RECT  9.56 104.895 11.54 104.965 ;
     RECT  11.08 16.695 11.61 16.765 ;
     RECT  11.46 42.035 11.65 42.525 ;
     RECT  9.88 47.495 11.65 48.265 ;
     RECT  11.08 53.235 11.65 53.725 ;
     RECT  11.27 57.435 11.65 60.445 ;
     RECT  9.88 68.775 11.65 68.985 ;
     RECT  11.65 42.035 11.84 49.385 ;
     RECT  11.84 40.915 12.03 49.385 ;
     RECT  11.65 53.235 12.03 61.845 ;
     RECT  12.03 40.915 12.22 61.845 ;
     RECT  12.03 65.835 12.22 65.905 ;
     RECT  11.65 68.775 12.22 69.685 ;
     RECT  10.01 26.915 12.41 26.985 ;
     RECT  12.22 40.915 12.41 70.245 ;
     RECT  12.41 40.915 12.6 71.785 ;
     RECT  11.46 32.095 12.79 33.705 ;
     RECT  11.46 36.855 12.79 38.045 ;
     RECT  12.6 40.915 12.98 71.925 ;
     RECT  13.55 23.695 13.74 23.765 ;
     RECT  12.41 26.915 13.93 28.525 ;
     RECT  12.79 32.095 13.93 38.045 ;
     RECT  13.74 23.695 14.12 24.045 ;
     RECT  13.55 83.755 14.31 83.825 ;
     RECT  13.93 26.915 14.5 38.045 ;
     RECT  12.98 40.915 14.5 75.985 ;
     RECT  14.12 22.715 14.69 24.045 ;
     RECT  14.5 26.915 14.69 75.985 ;
     RECT  10.21 79.135 14.69 79.205 ;
     RECT  14.31 83.755 14.69 84.525 ;
     RECT  14.69 21.595 15.22 75.985 ;
     RECT  14.69 79.135 15.22 84.525 ;
     RECT  5.2 88.375 15.22 90.545 ;
     RECT  15.22 16.31 15.68 90.545 ;
     RECT  11.12 0.035 20.02 0.105 ;
     RECT  11.54 104.755 20.02 104.965 ;
     RECT  15.68 16.975 20.345 90.545 ;
     RECT  20.345 16.835 20.68 90.545 ;
     RECT  20.02 0.035 21.12 8.63 ;
     RECT  20.02 94.97 21.12 98.23 ;
     RECT  20.02 103.37 21.12 104.965 ;
     RECT  20.68 16.835 23.81 87.185 ;
     RECT  20.68 90.335 23.81 90.545 ;
     RECT  23.81 16.835 25.22 90.545 ;
     RECT  25.22 16.31 25.68 90.545 ;
     RECT  21.12 0.035 30.02 0.105 ;
     RECT  25.14 10.395 30.02 10.465 ;
     RECT  30.02 0.035 31.12 10.465 ;
     RECT  30.02 93.57 31.12 99.63 ;
     RECT  25.68 17.115 31.41 90.545 ;
     RECT  31.41 16.975 35.22 90.545 ;
     RECT  35.22 16.31 35.68 90.545 ;
     RECT  31.12 10.395 39.58 10.465 ;
     RECT  35.68 16.975 39.96 90.545 ;
     RECT  31.12 0.035 40.02 0.105 ;
     RECT  39.58 9.135 40.02 10.465 ;
     RECT  21.12 104.755 40.02 104.965 ;
     RECT  40.02 0.035 41.12 10.465 ;
     RECT  40.02 94.97 41.12 98.23 ;
     RECT  40.02 103.37 41.12 104.965 ;
     RECT  39.96 16.835 45.22 90.545 ;
     RECT  45.22 16.31 45.68 90.545 ;
     RECT  41.12 0.035 50.02 0.385 ;
     RECT  41.12 9.135 50.02 10.465 ;
     RECT  41.12 95.795 50.02 95.865 ;
     RECT  50.02 0.035 51.12 10.465 ;
     RECT  50.02 93.57 51.12 99.63 ;
     RECT  45.68 16.835 51.81 90.545 ;
     RECT  51.12 9.135 54.635 10.465 ;
     RECT  51.12 95.795 55.16 95.865 ;
     RECT  51.81 17.115 55.22 90.545 ;
     RECT  55.22 16.31 55.68 90.545 ;
     RECT  55.68 16.975 58.58 19.705 ;
     RECT  55.68 23.835 58.58 90.545 ;
     RECT  58.58 16.975 58.84 90.545 ;
     RECT  51.12 0.035 60.02 0.385 ;
     RECT  54.635 9.135 60.02 10.325 ;
     RECT  55.16 94.535 60.02 95.865 ;
     RECT  41.12 104.755 60.02 104.965 ;
     RECT  60.02 0.035 61.12 10.325 ;
     RECT  60.02 94.535 61.12 98.23 ;
     RECT  60.02 103.37 61.12 104.965 ;
     RECT  58.84 17.255 64.09 90.545 ;
     RECT  64.09 17.115 65.22 90.545 ;
     RECT  65.22 16.31 65.87 90.545 ;
     RECT  65.87 16.31 67.26 85.925 ;
     RECT  67.26 15.295 68.72 85.925 ;
     RECT  61.12 9.135 69.265 10.325 ;
     RECT  68.72 16.975 69.41 85.925 ;
     RECT  69.41 16.975 69.6 86.065 ;
     RECT  65.87 89.495 69.6 90.545 ;
     RECT  69.265 9.135 69.78 10.465 ;
     RECT  61.12 0.035 70.02 0.385 ;
     RECT  69.78 9.135 70.02 10.605 ;
     RECT  61.12 94.535 70.02 95.865 ;
     RECT  69.6 16.975 70.24 90.545 ;
     RECT  70.02 0.035 71.12 10.605 ;
     RECT  70.02 93.57 71.12 99.63 ;
     RECT  61.12 104.755 71.95 104.965 ;
     RECT  70.24 17.115 73.4 90.545 ;
     RECT  71.12 9.135 73.535 10.605 ;
     RECT  73.4 16.975 75.22 90.545 ;
     RECT  75.22 16.31 75.68 90.545 ;
     RECT  75.68 16.975 78.41 67.165 ;
     RECT  75.68 70.175 79.67 87.325 ;
     RECT  75.68 90.335 79.67 90.545 ;
     RECT  71.12 0.035 80.02 0.385 ;
     RECT  73.535 9.135 80.02 10.465 ;
     RECT  71.12 94.535 80.02 95.865 ;
     RECT  71.95 104.895 80.02 104.965 ;
     RECT  78.41 17.115 80.22 67.165 ;
     RECT  79.67 70.175 80.22 90.545 ;
     RECT  80.22 17.115 80.68 90.545 ;
     RECT  80.68 75.775 80.69 90.545 ;
     RECT  80.02 0.035 81.12 10.465 ;
     RECT  80.02 94.535 81.12 98.23 ;
     RECT  80.02 103.37 81.12 104.965 ;
     RECT  80.68 17.115 81.26 50.645 ;
     RECT  81.26 20.755 81.64 50.645 ;
     RECT  81.26 17.115 81.76 17.605 ;
     RECT  80.69 75.775 81.83 79.765 ;
     RECT  80.68 53.935 82.21 60.585 ;
     RECT  81.83 75.775 82.21 78.645 ;
     RECT  81.64 20.755 82.4 50.505 ;
     RECT  82.4 21.315 82.59 36.085 ;
     RECT  82.21 54.915 82.59 60.585 ;
     RECT  80.69 82.775 82.59 90.545 ;
     RECT  82.59 32.795 82.78 36.085 ;
     RECT  82.59 54.915 82.78 59.185 ;
     RECT  82.59 82.775 82.78 82.985 ;
     RECT  81.76 16.975 82.97 17.605 ;
     RECT  82.4 38.955 82.97 50.505 ;
     RECT  82.78 56.175 82.97 59.185 ;
     RECT  82.21 78.015 82.97 78.645 ;
     RECT  82.59 85.855 82.97 90.545 ;
     RECT  82.97 17.535 83.16 17.605 ;
     RECT  82.78 33.635 83.16 36.085 ;
     RECT  82.97 85.855 83.16 87.045 ;
     RECT  82.59 21.315 83.35 29.925 ;
     RECT  82.97 44.555 83.35 50.505 ;
     RECT  83.16 85.855 83.35 85.925 ;
     RECT  83.16 35.315 83.54 36.085 ;
     RECT  82.97 38.955 83.54 40.985 ;
     RECT  83.35 44.555 83.54 48.125 ;
     RECT  80.68 66.955 83.54 68.565 ;
     RECT  82.78 82.775 83.54 82.845 ;
     RECT  83.35 24.115 83.73 29.925 ;
     RECT  83.54 46.655 83.73 48.125 ;
     RECT  83.54 39.235 83.92 40.985 ;
     RECT  83.73 46.655 83.92 47.985 ;
     RECT  83.54 35.875 83.93 36.085 ;
     RECT  83.73 29.855 84.11 29.925 ;
     RECT  83.92 40.915 84.11 40.985 ;
     RECT  82.97 89.915 84.11 90.545 ;
     RECT  83.73 24.115 84.3 25.445 ;
     RECT  82.97 57.295 84.68 59.185 ;
     RECT  83.54 66.955 84.88 68.005 ;
     RECT  82.97 78.435 84.88 78.645 ;
     RECT  81.12 0.035 84.9 0.385 ;
     RECT  84.88 78.435 84.97 78.505 ;
     RECT  81.12 104.895 85.18 104.965 ;
     RECT  84.9 0.035 85.25 0.525 ;
     RECT  84.3 25.375 85.25 25.445 ;
     RECT  83.93 36.015 85.25 36.085 ;
     RECT  81.12 9.135 85.46 10.465 ;
     RECT  83.92 46.655 85.53 46.725 ;
     RECT  84.88 67.935 85.53 68.005 ;
     RECT  85.25 0.315 85.81 0.525 ;
     RECT  84.68 57.295 85.81 57.365 ;
     RECT  85.46 8.995 88.165 10.465 ;
     RECT  85.81 0.455 90.02 0.525 ;
     RECT  88.165 8.995 90.02 10.605 ;
     RECT  84.11 89.915 90.02 90.405 ;
     RECT  81.12 94.535 90.02 95.865 ;
     RECT  90.02 54.37 90.69 57.63 ;
     RECT  90.02 0.455 91.12 10.605 ;
     RECT  90.02 15.17 91.12 18.43 ;
     RECT  90.02 23.57 91.12 29.63 ;
     RECT  90.02 34.77 91.12 38.03 ;
     RECT  90.02 43.17 91.12 49.23 ;
     RECT  90.02 62.77 91.12 68.83 ;
     RECT  90.02 73.97 91.12 80.03 ;
     RECT  90.02 85.17 91.12 90.405 ;
     RECT  90.02 93.57 91.12 99.63 ;
     RECT  91.12 8.995 91.69 10.605 ;
     RECT  90.69 54.37 91.83 58.205 ;
     RECT  91.12 62.77 91.83 68.005 ;
     RECT  91.83 54.37 92.97 68.005 ;
     RECT  92.97 54.215 93.73 68.005 ;
     RECT  93.73 52.395 94.87 68.005 ;
     RECT  91.12 0.455 95.5 0.525 ;
     RECT  91.69 8.995 95.5 10.465 ;
     RECT  94.87 47.355 95.5 47.425 ;
     RECT  94.87 51.975 95.5 68.005 ;
     RECT  91.12 90.335 95.5 90.405 ;
     RECT  91.12 94.535 95.5 95.865 ;
     RECT  85.18 104.755 95.5 104.965 ;
     RECT  95.5 0.455 96.2 104.965 ;
     RECT  96.2 0.455 98.665 0.525 ;
     RECT  96.2 90.335 99.24 90.405 ;
     RECT  96.2 94.535 99.46 95.865 ;
     RECT  98.665 0.175 100.02 0.525 ;
     RECT  96.2 8.995 100.02 10.465 ;
     RECT  99.24 22.295 100.02 22.365 ;
     RECT  96.2 34.615 100.02 68.285 ;
     RECT  99.46 73.535 100.02 73.605 ;
     RECT  99.24 90.335 100.02 90.545 ;
     RECT  99.46 94.535 100.02 96.005 ;
     RECT  96.2 104.755 100.02 104.965 ;
     RECT  100.02 73.535 100.26 78.63 ;
     RECT  100.02 33.37 100.64 68.285 ;
     RECT  100.02 0.175 101.12 10.465 ;
     RECT  100.02 13.77 101.12 28.23 ;
     RECT  100.64 33.37 101.12 59.03 ;
     RECT  100.26 75.37 101.12 78.63 ;
     RECT  100.02 83.77 101.12 90.545 ;
     RECT  100.02 94.535 101.12 98.23 ;
     RECT  100.02 103.37 101.12 104.965 ;
     RECT  101.12 34.615 101.21 58.205 ;
     RECT  100.64 61.915 101.21 68.145 ;
     RECT  101.21 34.615 101.49 46.865 ;
     RECT  101.21 61.915 101.59 65.345 ;
     RECT  101.49 39.935 101.78 46.865 ;
     RECT  101.49 34.615 101.97 37.065 ;
     RECT  101.78 39.935 101.97 42.525 ;
     RECT  101.78 45.535 101.97 46.865 ;
     RECT  101.21 50.155 101.97 58.205 ;
     RECT  101.59 65.275 101.97 65.345 ;
     RECT  101.97 50.155 102.16 51.765 ;
     RECT  101.97 56.175 102.35 58.205 ;
     RECT  102.16 50.295 102.54 51.765 ;
     RECT  102.35 56.595 102.54 58.205 ;
     RECT  102.54 57.015 102.73 58.205 ;
     RECT  101.12 90.335 104.56 90.545 ;
     RECT  101.12 94.535 104.56 96.005 ;
     RECT  104.56 90.335 104.85 96.005 ;
     RECT  101.97 34.615 104.88 34.685 ;
     RECT  104.78 81.095 104.88 81.165 ;
     RECT  104.37 68.775 105.51 68.845 ;
     RECT  105.51 67.655 105.7 68.845 ;
     RECT  101.12 22.295 105.89 22.365 ;
     RECT  105.7 29.715 105.89 29.785 ;
     RECT  102.73 57.015 105.89 57.925 ;
     RECT  105.51 62.475 105.89 62.545 ;
     RECT  105.51 53.655 106.08 53.725 ;
     RECT  105.89 57.015 106.08 58.345 ;
     RECT  105.89 61.215 106.08 62.545 ;
     RECT  105.7 66.675 106.08 68.845 ;
     RECT  105.89 85.995 106.08 86.065 ;
     RECT  105.89 22.295 106.27 24.745 ;
     RECT  105.89 27.615 106.27 29.785 ;
     RECT  101.97 45.535 106.27 45.605 ;
     RECT  106.08 53.655 106.27 68.845 ;
     RECT  106.27 21.875 106.46 29.785 ;
     RECT  104.88 33.775 106.46 34.685 ;
     RECT  106.27 53.655 106.46 71.085 ;
     RECT  104.88 80.255 106.46 81.165 ;
     RECT  106.08 85.995 106.46 87.885 ;
     RECT  106.27 45.535 106.84 46.305 ;
     RECT  106.65 49.875 106.84 49.945 ;
     RECT  106.46 52.815 106.84 71.085 ;
     RECT  104.85 92.015 106.91 96.005 ;
     RECT  106.84 38.955 107.03 39.025 ;
     RECT  106.84 45.535 107.03 49.945 ;
     RECT  106.84 52.815 107.03 73.465 ;
     RECT  106.46 18.655 107.22 34.685 ;
     RECT  107.03 38.675 107.22 40.145 ;
     RECT  107.03 45.535 107.22 73.605 ;
     RECT  107.22 18.655 107.6 73.605 ;
     RECT  106.46 80.255 107.79 87.885 ;
     RECT  107.6 17.815 108.36 73.605 ;
     RECT  107.79 77.595 108.36 87.885 ;
     RECT  101.12 0.175 110.02 0.245 ;
     RECT  101.12 8.995 110.02 10.465 ;
     RECT  108.36 17.815 110.07 87.885 ;
     RECT  110.02 0.175 110.22 10.465 ;
     RECT  107.22 13.755 110.22 13.825 ;
     RECT  110.07 17.815 110.22 89.145 ;
     RECT  106.91 94.535 110.22 96.005 ;
     RECT  110.22 0.175 110.68 96.005 ;
     RECT  110.68 0.175 111.12 10.465 ;
     RECT  110.02 99.17 111.12 99.63 ;
     RECT  111.12 8.995 114.63 10.465 ;
     RECT  110.68 13.615 114.63 89.705 ;
     RECT  114.63 8.995 115.22 89.705 ;
     RECT  110.68 94.535 115.22 96.005 ;
     RECT  115.22 8.995 115.68 96.005 ;
     RECT  115.68 8.995 119.19 91.665 ;
     RECT  115.68 94.535 119.19 96.005 ;
     RECT  111.12 0.175 120.02 0.245 ;
     RECT  119.19 8.995 120.02 96.005 ;
     RECT  101.12 104.755 120.02 104.965 ;
     RECT  120.02 0.175 121.12 5.83 ;
     RECT  120.02 8.995 121.12 98.23 ;
     RECT  120.02 103.37 121.12 104.965 ;
     RECT  121.12 8.995 125.91 96.005 ;
     RECT  121.12 0.175 127.81 0.245 ;
     RECT  125.91 8.995 130.02 91.665 ;
     RECT  130.02 1.17 130.22 91.665 ;
     RECT  125.91 94.535 130.22 96.005 ;
     RECT  130.22 1.17 130.68 96.005 ;
     RECT  130.68 1.17 131.12 76.125 ;
     RECT  130.02 99.17 131.12 99.63 ;
     RECT  131.12 8.995 134.2 76.125 ;
     RECT  134.2 8.995 134.77 76.405 ;
     RECT  134.77 8.995 135.22 76.545 ;
     RECT  130.68 80.675 135.22 90.405 ;
     RECT  130.68 94.535 135.22 96.005 ;
     RECT  135.22 8.995 135.68 96.005 ;
     RECT  135.68 8.995 139.52 15.785 ;
     RECT  135.68 18.655 139.52 89.285 ;
     RECT  135.68 92.855 140.02 96.005 ;
     RECT  121.12 104.755 140.02 104.965 ;
     RECT  139.52 8.995 140.22 89.285 ;
     RECT  140.02 92.855 140.22 98.23 ;
     RECT  140.02 2.57 141.12 5.83 ;
     RECT  140.22 8.995 141.12 98.23 ;
     RECT  140.02 103.37 141.12 104.965 ;
     RECT  141.12 8.995 146.81 96.005 ;
     RECT  146.81 67.935 149.4 96.005 ;
     RECT  149.4 67.935 149.74 98.805 ;
     RECT  149.74 67.655 149.78 98.805 ;
     RECT  146.81 8.995 150.02 63.945 ;
     RECT  149.78 67.515 150.02 98.805 ;
     RECT  150.02 1.17 150.22 63.945 ;
     RECT  150.02 67.515 150.22 99.63 ;
     RECT  150.22 1.17 151.12 99.63 ;
     RECT  141.12 104.755 156.69 104.965 ;
     RECT  156.69 104.895 160.02 104.965 ;
     RECT  160.02 2.57 161.12 5.83 ;
     RECT  160.02 103.37 161.12 104.965 ;
     RECT  151.12 8.995 170.02 98.805 ;
     RECT  170.02 1.17 171.12 99.63 ;
     RECT  171.12 8.995 172.08 98.805 ;
     RECT  172.08 8.995 175.22 10.465 ;
     RECT  172.08 13.335 175.22 98.805 ;
     RECT  175.22 8.995 175.68 98.805 ;
     RECT  175.68 8.995 179.04 10.465 ;
     RECT  175.68 13.335 179.04 92.085 ;
     RECT  179.04 8.995 179.42 92.085 ;
     RECT  175.68 95.935 179.42 98.805 ;
     RECT  161.12 104.895 180.02 104.965 ;
     RECT  179.42 8.995 181.01 98.805 ;
     RECT  180.02 2.57 181.12 5.83 ;
     RECT  180.02 103.37 181.12 104.965 ;
     RECT  181.01 92.015 181.58 98.805 ;
     RECT  181.01 8.995 185.22 89.145 ;
     RECT  181.58 92.015 185.22 92.225 ;
     RECT  181.58 95.935 185.22 98.805 ;
     RECT  185.22 8.995 185.68 98.805 ;
     RECT  185.68 21.875 185.95 89.145 ;
     RECT  185.95 30.275 186.52 89.145 ;
     RECT  186.52 30.275 186.71 89.005 ;
     RECT  181.12 104.895 186.865 104.965 ;
     RECT  186.71 30.275 186.9 46.585 ;
     RECT  186.865 104.755 186.935 104.965 ;
     RECT  186.71 49.735 187.09 89.005 ;
     RECT  186.9 30.275 187.28 45.605 ;
     RECT  185.68 14.315 187.47 18.725 ;
     RECT  187.09 50.575 187.47 89.005 ;
     RECT  185.95 21.875 187.66 26.005 ;
     RECT  187.28 36.435 187.66 45.605 ;
     RECT  187.47 50.575 187.66 56.805 ;
     RECT  187.66 25.795 187.85 26.005 ;
     RECT  187.28 30.275 187.85 33.145 ;
     RECT  187.66 36.855 187.85 45.605 ;
     RECT  187.66 52.535 187.85 56.805 ;
     RECT  187.47 61.075 187.85 79.345 ;
     RECT  187.85 45.535 188.04 45.605 ;
     RECT  187.85 63.315 188.04 79.345 ;
     RECT  187.47 83.055 188.04 89.005 ;
     RECT  187.47 16.275 188.23 18.725 ;
     RECT  187.66 21.875 188.23 21.945 ;
     RECT  187.85 30.275 188.23 32.165 ;
     RECT  187.85 56.735 188.23 56.805 ;
     RECT  188.04 63.315 188.23 78.225 ;
     RECT  187.85 36.855 188.42 41.965 ;
     RECT  188.23 73.395 188.42 78.225 ;
     RECT  188.42 74.935 188.61 78.225 ;
     RECT  188.04 83.055 188.61 84.805 ;
     RECT  188.61 74.935 188.8 77.945 ;
     RECT  187.85 25.795 188.99 25.865 ;
     RECT  188.23 63.315 188.99 68.565 ;
     RECT  188.61 83.055 188.99 83.125 ;
     RECT  188.42 36.855 189.37 36.925 ;
     RECT  185.68 95.935 189.37 98.805 ;
     RECT  188.99 63.875 189.56 66.045 ;
     RECT  189.37 98.735 189.69 98.805 ;
     RECT  188.23 30.275 189.81 30.485 ;
     RECT  188.23 17.815 189.88 18.725 ;
     RECT  189.81 29.575 189.88 30.485 ;
     RECT  188.42 41.755 189.88 41.965 ;
     RECT  187.85 52.535 189.88 53.445 ;
     RECT  189.56 65.135 189.88 66.045 ;
     RECT  188.8 76.615 189.88 77.525 ;
     RECT  188.04 87.675 189.88 89.005 ;
     RECT  189.88 29.575 189.94 29.645 ;
     RECT  185.68 8.995 189.97 10.465 ;
     RECT  189.88 52.535 189.97 52.605 ;
     RECT  189.88 65.975 189.97 66.045 ;
     RECT  190.02 1.17 191.12 7.23 ;
     RECT  190.02 99.17 191.12 99.63 ;
     RECT  189.97 10.395 195.5 10.465 ;
     RECT  186.935 104.755 195.5 104.825 ;
     RECT  195.5 1.33 195.64 104.825 ;
     RECT  195.64 2.73 196.2 104.825 ;
     RECT  196.2 104.755 198.87 104.825 ;
     RECT  196.2 10.395 199.965 10.465 ;
     RECT  199.75 41.755 199.965 41.825 ;
     RECT  199.75 72.835 199.965 72.905 ;
    LAYER metal4 ;
     RECT  85.705 0.28 85.845 0.42 ;
     RECT  84.865 0.42 85.845 1.17 ;
     RECT  10.02 1.17 11.12 1.33 ;
     RECT  84.865 1.17 91.12 1.33 ;
     RECT  190.02 1.17 191.12 1.33 ;
     RECT  84.865 1.33 95.64 2.57 ;
     RECT  190.02 1.33 195.64 2.73 ;
     RECT  120.02 2.57 121.12 5.83 ;
     RECT  140.02 2.57 141.12 5.83 ;
     RECT  160.02 2.57 161.12 5.83 ;
     RECT  180.02 2.57 181.12 5.83 ;
     RECT  110.02 1.17 111.12 7.23 ;
     RECT  20.02 2.57 21.12 8.63 ;
     RECT  40.02 2.57 41.12 8.63 ;
     RECT  60.02 2.57 61.12 8.63 ;
     RECT  80.02 2.57 101.12 8.63 ;
     RECT  190.02 2.73 196.2 8.96 ;
     RECT  4.5 1.33 11.12 10.03 ;
     RECT  30.02 1.17 31.12 10.03 ;
     RECT  50.02 1.17 51.12 10.03 ;
     RECT  70.02 1.17 71.12 10.03 ;
     RECT  170.02 1.17 171.12 12.04 ;
     RECT  110.22 7.23 111.12 12.67 ;
     RECT  120.22 5.83 120.68 12.67 ;
     RECT  130.02 1.17 131.12 12.67 ;
     RECT  140.22 5.83 140.68 12.67 ;
     RECT  150.02 1.17 151.12 12.67 ;
     RECT  160.22 5.83 160.68 12.67 ;
     RECT  169.585 12.04 171.12 12.67 ;
     RECT  180.22 5.83 180.68 12.67 ;
     RECT  189.865 8.96 196.2 12.67 ;
     RECT  4.5 10.03 5.2 15.68 ;
     RECT  0.585 15.68 5.2 15.96 ;
     RECT  67.225 15.26 67.365 16.31 ;
     RECT  15.22 16.31 15.68 16.66 ;
     RECT  45.22 16.31 45.68 16.94 ;
     RECT  11.505 16.66 15.68 17.71 ;
     RECT  25.22 16.31 25.68 17.71 ;
     RECT  35.22 16.31 35.68 17.71 ;
     RECT  44.905 16.94 45.68 17.71 ;
     RECT  55.22 16.31 55.68 17.71 ;
     RECT  65.22 16.31 67.365 17.71 ;
     RECT  75.22 16.31 75.68 17.71 ;
     RECT  84.865 8.63 101.12 17.71 ;
     RECT  110.22 12.67 196.2 17.78 ;
     RECT  108.825 17.78 196.2 24.78 ;
     RECT  108.265 24.78 196.2 25.62 ;
     RECT  106.865 25.62 196.2 30.38 ;
     RECT  11.505 17.71 101.12 39.62 ;
     RECT  11.505 39.62 101.245 39.76 ;
     RECT  107.145 30.38 196.2 39.76 ;
     RECT  11.505 39.76 196.2 40.18 ;
     RECT  107.425 40.18 196.2 44.38 ;
     RECT  110.22 44.38 196.2 52.64 ;
     RECT  11.505 40.18 101.805 53.9 ;
     RECT  110.22 52.64 189.725 57.68 ;
     RECT  0.025 15.96 5.2 58.1 ;
     RECT  11.505 53.9 101.12 58.1 ;
     RECT  108.545 57.68 189.725 64.96 ;
     RECT  107.705 64.96 189.725 65.94 ;
     RECT  195.5 52.64 196.2 65.94 ;
     RECT  0.025 58.1 101.12 67.43 ;
     RECT  107.705 65.94 196.2 71.54 ;
     RECT  0.025 67.43 99.565 75.37 ;
     RECT  0.025 75.37 101.12 81.06 ;
     RECT  109.665 71.54 196.2 81.06 ;
     RECT  0.025 81.06 196.2 87.85 ;
     RECT  0.025 87.85 15.68 89.25 ;
     RECT  25.22 87.85 25.68 89.25 ;
     RECT  35.22 87.85 35.68 89.25 ;
     RECT  45.22 87.85 45.68 89.25 ;
     RECT  55.22 87.85 55.68 89.25 ;
     RECT  65.22 87.85 65.68 89.25 ;
     RECT  73.745 87.85 75.68 89.25 ;
     RECT  73.745 89.25 73.885 89.74 ;
     RECT  85.145 87.85 196.2 90.44 ;
     RECT  110.22 90.44 196.2 92.61 ;
     RECT  115.22 92.61 125.68 94.01 ;
     RECT  135.22 92.61 145.68 94.01 ;
     RECT  155.22 92.61 165.68 94.01 ;
     RECT  175.22 92.61 196.2 94.01 ;
     RECT  0.025 89.25 12.205 94.5 ;
     RECT  189.305 94.01 196.2 94.78 ;
     RECT  85.145 90.44 101.12 94.97 ;
     RECT  4.5 94.5 12.205 95.9 ;
     RECT  189.585 94.78 196.2 98.84 ;
     RECT  4.5 95.9 11.645 99.63 ;
     RECT  30.02 93.57 31.12 99.63 ;
     RECT  50.02 93.57 51.12 99.63 ;
     RECT  70.02 93.57 71.12 99.63 ;
     RECT  80.02 94.97 101.12 99.63 ;
     RECT  110.02 99.17 111.12 99.63 ;
     RECT  130.02 99.17 131.12 99.63 ;
     RECT  150.02 99.17 151.12 99.63 ;
     RECT  170.02 99.17 171.12 99.63 ;
     RECT  190.02 98.84 196.2 99.63 ;
     RECT  4.5 99.63 5.2 102.27 ;
     RECT  95.5 99.63 101.12 102.27 ;
     RECT  195.5 99.63 196.2 102.27 ;
     RECT  5.06 102.27 5.2 103.67 ;
     RECT  96.06 102.27 101.12 103.67 ;
     RECT  196.06 102.27 196.2 103.67 ;
     RECT  20.02 94.97 21.12 103.83 ;
     RECT  40.02 94.97 41.12 103.83 ;
     RECT  60.02 94.97 61.12 103.83 ;
     RECT  80.02 99.63 85.285 103.83 ;
     RECT  100.02 103.67 101.12 103.83 ;
     RECT  120.02 94.01 121.12 103.83 ;
     RECT  140.02 94.01 141.12 103.83 ;
     RECT  160.02 94.01 161.12 103.83 ;
     RECT  180.02 94.01 181.12 103.83 ;
     RECT  11.505 99.63 11.645 104.86 ;
     RECT  85.145 103.83 85.285 104.86 ;
    LAYER metal5 ;
     RECT  0.025 15.96 0.585 16.1 ;
     RECT  0.585 15.68 4.5 16.1 ;
     RECT  4.5 1.33 5.06 102.27 ;
     RECT  5.06 1.33 5.2 103.67 ;
     RECT  5.2 1.33 10.05 10.02 ;
     RECT  10.05 1.18 11.09 10.02 ;
     RECT  5.2 89.6 11.09 99.62 ;
     RECT  5.2 15.68 15.23 16.1 ;
     RECT  11.09 89.6 15.23 90.02 ;
     RECT  15.23 15.68 20.05 90.02 ;
     RECT  11.09 95.76 20.05 95.9 ;
     RECT  20.05 2.58 21.09 8.62 ;
     RECT  20.05 15.68 21.09 103.82 ;
     RECT  21.09 15.68 30.05 90.02 ;
     RECT  21.09 95.76 30.05 95.9 ;
     RECT  30.05 1.18 31.09 10.02 ;
     RECT  30.05 15.68 31.09 99.62 ;
     RECT  31.09 15.68 40.05 90.02 ;
     RECT  31.09 95.76 40.05 95.9 ;
     RECT  40.05 2.58 41.09 8.62 ;
     RECT  40.05 15.68 41.09 103.82 ;
     RECT  41.09 15.68 50.05 90.02 ;
     RECT  41.09 95.76 50.05 95.9 ;
     RECT  50.05 1.18 51.09 10.02 ;
     RECT  50.05 15.68 51.09 99.62 ;
     RECT  51.09 15.68 60.05 90.02 ;
     RECT  51.09 95.76 60.05 95.9 ;
     RECT  60.05 2.58 61.09 8.62 ;
     RECT  60.05 15.68 61.09 103.82 ;
     RECT  61.09 15.68 67.365 90.02 ;
     RECT  67.365 15.96 70.05 90.02 ;
     RECT  61.09 95.76 70.05 95.9 ;
     RECT  70.05 1.18 71.09 10.02 ;
     RECT  70.05 15.96 71.09 99.62 ;
     RECT  71.09 15.96 74.645 90.02 ;
     RECT  74.645 16.31 75.67 90.02 ;
     RECT  75.67 17.71 80.05 90.02 ;
     RECT  71.09 95.76 80.05 95.9 ;
     RECT  80.05 17.71 80.67 103.82 ;
     RECT  80.67 89.88 80.805 103.82 ;
     RECT  80.05 2.58 81.09 8.62 ;
     RECT  80.805 94.64 81.09 103.82 ;
     RECT  85.145 10.64 90.05 10.78 ;
     RECT  81.09 94.64 90.05 95.9 ;
     RECT  90.05 1.18 91.09 99.62 ;
     RECT  91.09 1.33 95.5 99.62 ;
     RECT  95.5 1.33 95.64 102.27 ;
     RECT  95.64 2.58 96.06 102.27 ;
     RECT  96.06 2.58 96.2 103.67 ;
     RECT  96.2 75.38 100.05 103.67 ;
     RECT  96.2 2.58 101.09 67.42 ;
     RECT  100.05 75.38 101.09 103.82 ;
     RECT  101.09 94.36 101.525 95.9 ;
     RECT  101.09 10.64 110.05 10.78 ;
     RECT  101.525 94.64 110.05 95.9 ;
     RECT  110.05 1.18 110.23 10.78 ;
     RECT  110.05 94.64 110.23 99.62 ;
     RECT  110.23 1.18 111.09 99.62 ;
     RECT  111.09 10.64 120.05 95.9 ;
     RECT  120.05 2.58 121.09 103.82 ;
     RECT  121.09 10.64 130.05 95.9 ;
     RECT  130.05 1.18 131.09 99.62 ;
     RECT  131.09 10.64 140.05 95.9 ;
     RECT  140.05 2.58 141.09 103.82 ;
     RECT  141.09 10.64 150.05 95.9 ;
     RECT  150.05 1.18 151.09 99.62 ;
     RECT  151.09 10.64 160.05 95.9 ;
     RECT  160.05 2.58 161.09 103.82 ;
     RECT  161.09 10.64 170.05 95.9 ;
     RECT  170.05 1.18 171.09 99.62 ;
     RECT  171.09 12.67 180.05 95.9 ;
     RECT  180.05 2.58 180.23 5.82 ;
     RECT  180.05 12.67 180.23 103.82 ;
     RECT  180.23 2.58 180.67 103.82 ;
     RECT  180.67 2.58 181.09 5.82 ;
     RECT  180.67 12.67 181.09 103.82 ;
     RECT  181.09 12.67 185.67 95.9 ;
     RECT  185.67 94.64 189.445 95.9 ;
     RECT  189.445 95.76 190.05 95.9 ;
     RECT  190.05 1.18 191.09 7.22 ;
     RECT  191.09 1.33 195.5 7.22 ;
     RECT  190.05 95.76 195.5 99.62 ;
     RECT  195.5 1.33 195.64 102.27 ;
     RECT  195.64 2.73 196.06 102.27 ;
     RECT  196.06 2.73 196.2 103.67 ;
    LAYER metal6 ;
     RECT  4.43 0 5.27 1.18 ;
     RECT  95.43 0 96.27 1.18 ;
     RECT  195.43 0 196.27 1.18 ;
     RECT  90.05 1.18 96.27 2.58 ;
     RECT  110.05 1.18 111.09 7.22 ;
     RECT  190.05 1.18 196.27 7.22 ;
     RECT  20.05 2.58 21.09 8.62 ;
     RECT  40.05 2.58 41.09 8.62 ;
     RECT  60.05 2.58 61.09 8.62 ;
     RECT  80.05 2.58 81.09 8.62 ;
     RECT  110.17 7.22 111.09 9.94 ;
     RECT  120.05 2.58 121.09 9.94 ;
     RECT  130.05 1.18 131.09 9.94 ;
     RECT  140.05 2.58 141.09 9.94 ;
     RECT  150.05 1.18 151.09 9.94 ;
     RECT  160.05 2.58 161.09 9.94 ;
     RECT  170.05 1.18 171.09 9.94 ;
     RECT  180.05 2.58 181.09 9.94 ;
     RECT  4.43 1.18 11.09 10.02 ;
     RECT  30.05 1.18 31.09 14.98 ;
     RECT  50.05 1.18 51.09 14.98 ;
     RECT  70.05 1.18 71.09 14.98 ;
     RECT  90.05 2.58 101.09 67.42 ;
     RECT  90.05 67.42 96.27 75.38 ;
     RECT  15.17 14.98 80.73 89.98 ;
     RECT  4.43 10.02 5.27 93.58 ;
     RECT  110.17 9.94 185.73 94.94 ;
     RECT  80.05 89.98 80.73 94.98 ;
     RECT  110.17 94.94 111.09 99.18 ;
     RECT  195.43 7.22 196.27 99.18 ;
     RECT  4.43 93.58 11.09 99.62 ;
     RECT  30.05 89.98 31.09 99.62 ;
     RECT  50.05 89.98 51.09 99.62 ;
     RECT  70.05 89.98 71.09 99.62 ;
     RECT  90.05 75.38 101.09 99.62 ;
     RECT  110.05 99.18 111.09 99.62 ;
     RECT  130.05 94.94 131.09 99.62 ;
     RECT  150.05 94.94 151.09 99.62 ;
     RECT  170.05 94.94 171.09 99.62 ;
     RECT  190.05 99.18 196.27 99.62 ;
     RECT  20.05 89.98 21.09 103.82 ;
     RECT  40.05 89.98 41.09 103.82 ;
     RECT  60.05 89.98 61.09 103.82 ;
     RECT  80.05 94.98 81.09 103.82 ;
     RECT  95.43 99.62 101.09 103.82 ;
     RECT  120.05 94.94 121.09 103.82 ;
     RECT  140.05 94.94 141.09 103.82 ;
     RECT  160.05 94.94 161.09 103.82 ;
     RECT  180.05 94.94 181.09 103.82 ;
     RECT  4.43 99.62 5.27 105 ;
     RECT  95.43 103.82 96.27 105 ;
     RECT  195.43 99.62 196.27 105 ;
    LAYER metal7 ;
     RECT  0 10.8 10.07 102 ;
     RECT  10.07 1.2 11.07 102 ;
     RECT  11.07 2.6 20.07 102 ;
     RECT  20.07 2.6 21.07 103.8 ;
     RECT  21.07 2.6 30.07 102 ;
     RECT  30.07 1.2 31.07 102 ;
     RECT  31.07 2.6 40.07 102 ;
     RECT  40.07 2.6 41.07 103.8 ;
     RECT  41.07 2.6 50.07 102 ;
     RECT  50.07 1.2 51.07 102 ;
     RECT  51.07 2.6 60.07 102 ;
     RECT  60.07 2.6 61.07 103.8 ;
     RECT  61.07 2.6 70.07 102 ;
     RECT  70.07 1.2 71.07 102 ;
     RECT  71.07 2.6 80.07 102 ;
     RECT  80.07 2.6 81.07 103.8 ;
     RECT  81.07 2.6 90.07 102 ;
     RECT  90.07 1.2 91.07 102 ;
     RECT  91.07 2.6 100.07 102 ;
     RECT  100.07 2.6 101.07 103.8 ;
     RECT  101.07 2.6 110.07 102 ;
     RECT  110.07 1.2 111.07 102 ;
     RECT  111.07 2.6 120.07 102 ;
     RECT  120.07 2.6 121.07 103.8 ;
     RECT  121.07 2.6 130.07 102 ;
     RECT  130.07 1.2 131.07 102 ;
     RECT  131.07 2.6 140.07 102 ;
     RECT  140.07 2.6 141.07 103.8 ;
     RECT  141.07 2.6 150.07 102 ;
     RECT  150.07 1.2 151.07 102 ;
     RECT  151.07 2.6 160.07 102 ;
     RECT  160.07 2.6 161.07 103.8 ;
     RECT  161.07 2.6 170.07 102 ;
     RECT  170.07 1.2 171.07 102 ;
     RECT  171.07 2.6 180.07 102 ;
     RECT  180.07 2.6 181.07 103.8 ;
     RECT  181.07 2.6 190.07 102 ;
     RECT  190.07 1.2 191.07 102 ;
     RECT  191.07 10.8 200 102 ;
    LAYER metal8 ;
     RECT  9.97 0 191.17 105 ;
  END
END top
END LIBRARY
