VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

VIA via1_2_1120_340_1_3_300_300
  VIARULE Via1Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal1 via1 metal2 ;
  CUTSPACING 0.08 0.08 ;
  ENCLOSURE 0.035 0.05 0.035 0.035 ;
  ROWCOL 1 3 ;
END via1_2_1120_340_1_3_300_300

VIA via2_3_1120_340_1_3_320_320
  VIARULE Via2Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal2 via2 metal3 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.035 0.035 ;
  ROWCOL 1 3 ;
END via2_3_1120_340_1_3_320_320

VIA via3_4_1120_340_1_3_320_320
  VIARULE Via3Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal3 via3 metal4 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.035 0.035 ;
  ROWCOL 1 3 ;
END via3_4_1120_340_1_3_320_320

VIA via4_5_1120_340_1_2_600_600
  VIARULE Via4Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal4 via4 metal5 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0 0 ;
  ROWCOL 1 2 ;
END via4_5_1120_340_1_2_600_600

VIA via5_6_1120_340_1_2_600_600
  VIARULE Via5Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal5 via5 metal6 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0.06 0 ;
  ROWCOL 1 2 ;
END via5_6_1120_340_1_2_600_600

MACRO enfasi
  FOREIGN enfasi 0 0 ;
  CLASS BLOCK ;
  SIZE 85 BY 85 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  84.93 31.955 85 32.025 ;
    END
  END clk
  PIN q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 23.835 0.07 23.905 ;
    END
  END q[0]
  PIN q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  60.48 84.93 60.55 85 ;
    END
  END q[10]
  PIN q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  84.93 8.715 85 8.785 ;
    END
  END q[11]
  PIN q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  84.93 78.435 85 78.505 ;
    END
  END q[1]
  PIN q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  13.36 84.93 13.43 85 ;
    END
  END q[2]
  PIN q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 35.595 0.07 35.665 ;
    END
  END q[3]
  PIN q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  76.44 84.93 76.51 85 ;
    END
  END q[4]
  PIN q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 82.075 0.07 82.145 ;
    END
  END q[5]
  PIN q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  47.94 0 48.01 0.07 ;
    END
  END q[6]
  PIN q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.355 0.07 12.425 ;
    END
  END q[7]
  PIN q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  79.48 0 79.55 0.07 ;
    END
  END q[8]
  PIN q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  0.82 0 0.89 0.07 ;
    END
  END q[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  16.4 0 16.47 0.07 ;
    END
  END rst
  PIN z[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  28.94 84.93 29.01 85 ;
    END
  END z[0]
  PIN z[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  84.93 20.475 85 20.545 ;
    END
  END z[10]
  PIN z[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  31.98 0 32.05 0.07 ;
    END
  END z[1]
  PIN z[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  84.93 55.195 85 55.265 ;
    END
  END z[2]
  PIN z[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  84.93 66.675 85 66.745 ;
    END
  END z[3]
  PIN z[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 58.835 0.07 58.905 ;
    END
  END z[4]
  PIN z[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  44.9 84.93 44.97 85 ;
    END
  END z[5]
  PIN z[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  63.52 0 63.59 0.07 ;
    END
  END z[6]
  PIN z[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 47.075 0.07 47.145 ;
    END
  END z[7]
  PIN z[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 70.315 0.07 70.385 ;
    END
  END z[8]
  PIN z[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  84.93 43.435 85 43.505 ;
    END
  END z[9]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal6 ;
        RECT  75.29 84.86 75.85 85 ;
        RECT  75.29 0 75.85 0.14 ;
        RECT  65.29 84.86 65.85 85 ;
        RECT  65.29 0 65.85 0.14 ;
        RECT  55.29 84.86 55.85 85 ;
        RECT  55.29 0 55.85 0.14 ;
        RECT  45.29 84.86 45.85 85 ;
        RECT  45.29 0 45.85 0.14 ;
        RECT  35.29 84.86 35.85 85 ;
        RECT  35.29 0 35.85 0.14 ;
        RECT  25.29 84.86 25.85 85 ;
        RECT  25.29 0 25.85 0.14 ;
        RECT  15.29 84.86 15.85 85 ;
        RECT  15.29 0 15.85 0.14 ;
        RECT  5.29 84.86 5.85 85 ;
        RECT  5.29 0 5.85 0.14 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal6 ;
        RECT  80.29 84.86 80.85 85 ;
        RECT  80.29 0 80.85 0.14 ;
        RECT  70.29 84.86 70.85 85 ;
        RECT  70.29 0 70.85 0.14 ;
        RECT  60.29 84.86 60.85 85 ;
        RECT  60.29 0 60.85 0.14 ;
        RECT  50.29 84.86 50.85 85 ;
        RECT  50.29 0 50.85 0.14 ;
        RECT  40.29 84.86 40.85 85 ;
        RECT  40.29 0 40.85 0.14 ;
        RECT  30.29 84.86 30.85 85 ;
        RECT  30.29 0 30.85 0.14 ;
        RECT  20.29 84.86 20.85 85 ;
        RECT  20.29 0 20.85 0.14 ;
        RECT  10.29 84.86 10.85 85 ;
        RECT  10.29 0 10.85 0.14 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
     RECT  0.57 1.315 2.34 84.085 ;
     RECT  2.34 1.155 10.89 84.085 ;
     RECT  10.89 1.155 14.88 84.245 ;
     RECT  14.88 1.015 16.4 84.245 ;
     RECT  16.4 1.015 17.16 84.385 ;
     RECT  17.16 1.015 22.55 84.525 ;
     RECT  22.55 1.015 24.07 84.245 ;
     RECT  24.07 1.015 24.76 84.085 ;
     RECT  24.76 0.875 28.06 84.085 ;
     RECT  28.06 1.015 28.25 84.085 ;
     RECT  28.25 1.155 28.94 84.085 ;
     RECT  28.94 1.155 31.98 84.385 ;
     RECT  31.98 1.015 32.62 84.385 ;
     RECT  32.62 1.015 39.2 84.245 ;
     RECT  39.2 1.015 39.96 84.525 ;
     RECT  39.96 1.015 41.48 84.665 ;
     RECT  41.48 0.875 49.15 84.665 ;
     RECT  49.15 0.875 57.32 84.525 ;
     RECT  57.32 1.155 64.92 84.525 ;
     RECT  64.92 1.315 69.1 84.525 ;
     RECT  69.1 1.315 74.99 84.385 ;
     RECT  74.99 1.315 84.36 84.085 ;
     RECT  84.36 57.995 84.87 58.065 ;
    LAYER metal2 ;
     RECT  15.07 0 16.28 0.035 ;
     RECT  78.72 0 79.36 0.035 ;
     RECT  47.94 0.035 48.01 0.875 ;
     RECT  15.07 0.035 16.47 1.015 ;
     RECT  24.76 0.875 28.06 1.015 ;
     RECT  31.98 0.035 32.05 1.015 ;
     RECT  41.48 0.875 41.55 1.015 ;
     RECT  47.37 0.875 48.01 1.015 ;
     RECT  57.25 0.875 57.32 1.015 ;
     RECT  0.82 0.035 0.89 1.155 ;
     RECT  14.88 1.015 16.47 1.155 ;
     RECT  55.16 1.015 57.32 1.155 ;
     RECT  63.52 0.035 63.59 1.155 ;
     RECT  0.82 1.155 2.41 1.33 ;
     RECT  21.53 1.015 32.05 1.33 ;
     RECT  63.52 1.155 64.92 1.33 ;
     RECT  78.72 0.035 79.55 1.33 ;
     RECT  41.48 1.015 50.48 1.575 ;
     RECT  54.97 1.155 57.7 1.575 ;
     RECT  12.03 1.155 16.47 1.715 ;
     RECT  21.53 1.33 35.8 1.715 ;
     RECT  40.34 1.575 57.7 1.715 ;
     RECT  63.52 1.33 65.8 1.715 ;
     RECT  75.34 1.33 79.55 1.715 ;
     RECT  0.82 1.33 5.8 1.785 ;
     RECT  12.03 1.715 57.7 1.855 ;
     RECT  62.19 1.715 65.8 1.855 ;
     RECT  10.13 1.855 65.8 1.995 ;
     RECT  75.34 1.715 79.74 1.995 ;
     RECT  10.13 1.995 67.2 2.275 ;
     RECT  2.34 1.785 5.8 2.415 ;
     RECT  9.94 2.275 67.2 2.415 ;
     RECT  73.02 1.995 82.59 2.415 ;
     RECT  2.34 2.415 67.2 2.73 ;
     RECT  73.02 2.415 84.11 2.73 ;
     RECT  2.34 2.73 84.11 3.605 ;
     RECT  2.34 3.605 83.73 8.155 ;
     RECT  2.34 8.155 84.11 8.715 ;
     RECT  1.58 8.715 84.11 9.135 ;
     RECT  1.39 9.135 84.11 9.205 ;
     RECT  1.39 9.205 83.73 12.355 ;
     RECT  1.01 12.355 83.73 13.755 ;
     RECT  1.01 13.755 84.11 15.015 ;
     RECT  0.82 15.015 84.11 16.065 ;
     RECT  0.82 16.065 83.92 19.845 ;
     RECT  1.58 19.845 83.92 19.985 ;
     RECT  1.77 19.985 83.92 20.475 ;
     RECT  1.77 20.475 84.11 21.665 ;
     RECT  1.77 21.665 83.35 23.835 ;
     RECT  0.82 23.835 83.35 25.585 ;
     RECT  1.96 25.585 83.35 25.935 ;
     RECT  1.96 25.935 84.3 26.915 ;
     RECT  1.96 26.915 84.49 30.415 ;
     RECT  1.39 30.415 84.49 33.635 ;
     RECT  1.39 33.635 84.11 35.595 ;
     RECT  0.82 35.595 84.11 38.185 ;
     RECT  1.39 38.185 84.11 42.735 ;
     RECT  1.39 42.735 84.3 43.715 ;
     RECT  0.63 43.715 84.3 48.335 ;
     RECT  0.82 48.335 84.11 52.535 ;
     RECT  0.63 52.535 84.11 53.935 ;
     RECT  0.63 53.935 84.68 57.785 ;
     RECT  0.82 57.785 84.68 57.995 ;
     RECT  0.82 57.995 84.87 62.965 ;
     RECT  0.63 62.965 84.87 73.185 ;
     RECT  0.63 73.185 84.11 73.605 ;
     RECT  0.63 73.605 83.73 74.445 ;
     RECT  1.01 74.445 83.73 77.595 ;
     RECT  1.01 77.595 84.11 77.665 ;
     RECT  1.39 77.665 84.3 77.945 ;
     RECT  1.96 77.945 84.3 80.045 ;
     RECT  1.96 80.045 83.92 80.465 ;
     RECT  1.96 80.465 82.21 82.005 ;
     RECT  1.96 82.005 5.8 82.145 ;
     RECT  5.34 82.145 5.8 82.67 ;
     RECT  10.13 82.005 80.8 82.67 ;
     RECT  10.13 82.67 24.07 83.265 ;
     RECT  28.94 82.67 80.8 83.265 ;
     RECT  37.11 83.265 71 83.545 ;
     RECT  10.34 83.265 24.07 84.07 ;
     RECT  80.34 83.265 80.8 84.07 ;
     RECT  10.89 84.07 24.07 84.245 ;
     RECT  37.11 83.545 63.97 84.245 ;
     RECT  69.03 83.545 71 84.245 ;
     RECT  21.34 84.245 22.55 84.385 ;
     RECT  28.94 83.265 32.62 84.385 ;
     RECT  39.2 84.245 40.98 84.385 ;
     RECT  44.9 84.245 63.97 84.385 ;
     RECT  74.92 83.265 76.51 84.385 ;
     RECT  12.6 84.245 17.23 84.525 ;
     RECT  22.48 84.385 22.55 84.525 ;
     RECT  39.2 84.385 40.03 84.525 ;
     RECT  44.9 84.385 49.72 84.525 ;
     RECT  54.02 84.385 54.09 84.525 ;
     RECT  69.03 84.245 69.1 84.525 ;
     RECT  39.96 84.525 40.03 84.665 ;
     RECT  44.9 84.525 49.15 84.665 ;
     RECT  59.91 84.385 63.4 84.945 ;
     RECT  12.6 84.525 13.43 84.965 ;
     RECT  28.94 84.385 29.01 84.965 ;
     RECT  44.9 84.665 44.97 84.965 ;
     RECT  59.91 84.945 60.55 84.965 ;
     RECT  76.44 84.385 76.51 84.965 ;
     RECT  12.6 84.965 13.24 85 ;
     RECT  59.91 84.965 60.36 85 ;
    LAYER metal3 ;
     RECT  0.035 58.835 0.63 58.905 ;
     RECT  0.63 57.715 0.82 58.905 ;
     RECT  0.035 12.355 1.01 12.425 ;
     RECT  0.82 19.775 1.01 19.845 ;
     RECT  0.035 47.075 1.01 47.145 ;
     RECT  0.63 52.535 1.01 52.605 ;
     RECT  0.63 43.715 1.2 43.785 ;
     RECT  1.01 47.075 1.2 48.405 ;
     RECT  1.01 51.275 1.2 52.605 ;
     RECT  0.82 56.735 1.2 58.905 ;
     RECT  1.01 76.055 1.2 76.125 ;
     RECT  1.01 12.355 1.39 14.805 ;
     RECT  1.01 17.675 1.39 19.845 ;
     RECT  0.035 35.595 1.39 35.665 ;
     RECT  1.2 43.715 1.39 58.905 ;
     RECT  1.39 11.935 1.58 19.845 ;
     RECT  0.035 23.835 1.58 23.905 ;
     RECT  1.39 43.715 1.58 61.145 ;
     RECT  0.035 70.315 1.58 70.385 ;
     RECT  1.2 76.055 1.58 77.945 ;
     RECT  1.58 8.715 1.77 23.905 ;
     RECT  1.39 35.595 1.96 36.365 ;
     RECT  1.77 39.935 1.96 40.005 ;
     RECT  1.58 42.875 1.96 61.145 ;
     RECT  0.035 82.075 2.03 82.145 ;
     RECT  1.96 29.015 2.15 29.085 ;
     RECT  1.96 35.595 2.15 40.005 ;
     RECT  1.96 42.875 2.15 63.525 ;
     RECT  1.77 8.715 2.34 24.465 ;
     RECT  2.15 28.735 2.34 30.205 ;
     RECT  2.15 35.595 2.34 63.665 ;
     RECT  2.34 8.715 2.72 63.665 ;
     RECT  1.58 70.315 2.91 77.945 ;
     RECT  2.72 7.875 3.48 63.665 ;
     RECT  2.91 67.655 3.48 77.945 ;
     RECT  3.48 7.875 5.19 77.945 ;
     RECT  2.34 3.815 5.34 3.885 ;
     RECT  5.19 7.875 5.34 79.205 ;
     RECT  5.34 1.33 5.8 82.67 ;
     RECT  5.8 3.675 9.75 79.765 ;
     RECT  9.75 3.255 9.94 79.765 ;
     RECT  9.94 3.115 10.34 79.765 ;
     RECT  10.34 2.73 10.8 84.07 ;
     RECT  10.8 2.73 12.98 81.725 ;
     RECT  12.98 2.555 14.31 81.725 ;
     RECT  14.31 2.555 15.34 82.005 ;
     RECT  15.34 1.33 15.8 82.67 ;
     RECT  15.8 1.995 19.82 82.005 ;
     RECT  19.82 1.855 20.34 82.005 ;
     RECT  20.34 1.855 20.8 84.07 ;
     RECT  20.8 1.855 21.03 82.005 ;
     RECT  21.03 1.855 21.15 81.725 ;
     RECT  21.15 1.715 21.98 81.725 ;
     RECT  21.98 1.995 25.34 81.725 ;
     RECT  25.34 1.33 25.8 82.67 ;
     RECT  25.8 1.995 29.32 66.185 ;
     RECT  29.32 1.995 29.89 66.465 ;
     RECT  29.89 1.995 30.34 66.605 ;
     RECT  25.8 70.735 30.34 80.465 ;
     RECT  30.34 1.995 30.72 84.07 ;
     RECT  30.72 2.275 30.8 84.07 ;
     RECT  30.8 2.275 34.64 5.845 ;
     RECT  30.8 8.715 34.64 79.345 ;
     RECT  34.64 2.275 35.34 79.345 ;
     RECT  30.8 82.915 35.34 82.985 ;
     RECT  35.34 1.33 35.8 82.985 ;
     RECT  35.8 1.715 37.3 82.985 ;
     RECT  37.3 1.715 40.34 83.265 ;
     RECT  40.34 1.575 40.8 84.07 ;
     RECT  40.8 1.575 41.93 83.265 ;
     RECT  41.93 57.995 44.86 83.265 ;
     RECT  44.86 57.715 44.9 83.265 ;
     RECT  41.93 1.575 45.34 54.005 ;
     RECT  44.9 57.575 45.34 84.945 ;
     RECT  45.34 1.33 45.8 84.945 ;
     RECT  45.8 1.575 55.34 84.945 ;
     RECT  55.34 1.33 55.8 84.945 ;
     RECT  55.8 1.715 58.27 84.945 ;
     RECT  58.27 2.275 62.19 84.945 ;
     RECT  62.19 1.715 63.4 84.945 ;
     RECT  63.4 1.715 65.34 83.405 ;
     RECT  65.34 1.33 65.8 83.405 ;
     RECT  65.8 1.715 66.06 83.405 ;
     RECT  66.06 1.715 67.01 83.265 ;
     RECT  67.01 3.255 67.2 83.265 ;
     RECT  67.2 3.395 70.34 83.265 ;
     RECT  70.34 2.73 70.8 84.07 ;
     RECT  70.8 3.395 74.16 82.145 ;
     RECT  74.16 3.115 74.54 82.145 ;
     RECT  74.54 3.115 75.34 83.265 ;
     RECT  75.34 1.33 75.8 83.265 ;
     RECT  75.8 1.995 76.13 83.265 ;
     RECT  76.13 82.075 76.7 83.265 ;
     RECT  76.13 1.995 79.55 79.205 ;
     RECT  79.55 2.73 80.34 79.205 ;
     RECT  76.7 82.075 80.34 82.285 ;
     RECT  80.34 2.73 80.8 84.07 ;
     RECT  80.8 11.935 81.07 79.205 ;
     RECT  81.07 20.335 81.64 79.205 ;
     RECT  81.64 20.335 81.83 79.065 ;
     RECT  81.83 20.335 82.02 36.645 ;
     RECT  81.83 39.795 82.21 79.065 ;
     RECT  82.02 20.335 82.4 35.665 ;
     RECT  80.8 4.375 82.59 8.785 ;
     RECT  82.4 20.335 82.59 23.205 ;
     RECT  82.21 40.635 82.59 79.065 ;
     RECT  81.07 11.935 82.78 16.065 ;
     RECT  82.4 26.495 82.78 35.665 ;
     RECT  82.59 40.635 82.78 46.865 ;
     RECT  82.78 15.855 82.97 16.065 ;
     RECT  82.59 20.475 82.97 23.205 ;
     RECT  82.78 26.915 82.97 35.665 ;
     RECT  82.78 42.735 82.97 46.865 ;
     RECT  82.59 51.135 82.97 69.405 ;
     RECT  82.97 35.595 83.16 35.665 ;
     RECT  82.97 53.375 83.16 69.405 ;
     RECT  82.59 73.115 83.16 79.065 ;
     RECT  82.59 6.335 83.35 8.785 ;
     RECT  82.78 11.935 83.35 12.005 ;
     RECT  82.97 20.475 83.35 22.225 ;
     RECT  82.97 46.795 83.35 46.865 ;
     RECT  83.16 53.375 83.35 68.285 ;
     RECT  83.16 77.735 83.35 79.065 ;
     RECT  82.97 26.915 83.54 32.025 ;
     RECT  82.97 42.735 83.54 43.505 ;
     RECT  83.35 63.455 83.54 68.285 ;
     RECT  83.35 53.375 83.73 58.625 ;
     RECT  83.54 64.995 83.73 68.285 ;
     RECT  83.16 73.115 83.73 74.865 ;
     RECT  83.73 64.995 83.92 68.005 ;
     RECT  82.97 15.855 84.11 15.925 ;
     RECT  83.73 53.375 84.11 55.265 ;
     RECT  83.73 58.555 84.11 58.625 ;
     RECT  83.73 73.115 84.11 73.185 ;
     RECT  83.54 26.915 84.49 26.985 ;
     RECT  84.11 53.935 84.68 55.265 ;
     RECT  83.35 8.715 84.965 8.785 ;
     RECT  83.35 20.475 84.965 20.545 ;
     RECT  83.54 31.955 84.965 32.025 ;
     RECT  83.54 43.435 84.965 43.505 ;
     RECT  84.68 55.195 84.965 55.265 ;
     RECT  83.92 66.675 84.965 66.745 ;
     RECT  83.35 77.735 84.965 78.505 ;
     RECT  84.965 77.735 85 78.365 ;
    LAYER metal4 ;
     RECT  65.34 1.33 65.8 2.1 ;
     RECT  5.34 1.33 5.8 2.73 ;
     RECT  15.34 1.33 15.8 2.73 ;
     RECT  25.34 1.33 25.8 2.73 ;
     RECT  35.34 1.33 35.8 2.73 ;
     RECT  45.34 1.33 45.8 2.73 ;
     RECT  55.34 1.33 55.8 2.73 ;
     RECT  64.705 2.1 65.8 2.73 ;
     RECT  75.34 1.33 75.8 2.73 ;
     RECT  5.34 2.73 80.8 7.84 ;
     RECT  3.945 7.84 80.8 14.84 ;
     RECT  3.385 14.84 80.8 15.68 ;
     RECT  1.985 15.68 80.8 20.44 ;
     RECT  2.265 20.44 80.8 30.24 ;
     RECT  2.545 30.24 80.8 33.18 ;
     RECT  2.545 33.18 81.925 34.44 ;
     RECT  5.34 34.44 81.925 47.74 ;
     RECT  3.665 47.74 81.925 52.5 ;
     RECT  3.665 52.5 81.365 52.92 ;
     RECT  3.665 52.92 80.8 55.02 ;
     RECT  2.825 55.02 80.8 61.6 ;
     RECT  4.785 61.6 80.8 72.94 ;
     RECT  5.34 72.94 80.8 82.67 ;
     RECT  10.34 82.67 10.8 84.07 ;
     RECT  20.34 82.67 20.8 84.07 ;
     RECT  30.34 82.67 30.8 84.07 ;
     RECT  40.34 82.67 40.8 84.07 ;
     RECT  50.34 82.67 50.8 84.07 ;
     RECT  60.34 82.67 60.8 84.07 ;
     RECT  70.34 82.67 70.8 84.07 ;
     RECT  80.34 82.67 80.8 84.07 ;
    LAYER metal5 ;
     RECT  5.35 1.33 5.79 82.67 ;
     RECT  5.79 2.73 10.35 82.67 ;
     RECT  10.35 2.73 10.79 84.07 ;
     RECT  10.79 2.73 15.35 82.67 ;
     RECT  15.35 1.33 15.79 82.67 ;
     RECT  15.79 2.73 20.35 82.67 ;
     RECT  20.35 2.73 20.79 84.07 ;
     RECT  20.79 2.73 25.35 82.67 ;
     RECT  25.35 1.33 25.79 82.67 ;
     RECT  25.79 2.73 30.35 82.67 ;
     RECT  30.35 2.73 30.79 84.07 ;
     RECT  30.79 2.73 35.35 82.67 ;
     RECT  35.35 1.33 35.79 82.67 ;
     RECT  35.79 2.73 40.35 82.67 ;
     RECT  40.35 2.73 40.79 84.07 ;
     RECT  40.79 2.73 45.35 82.67 ;
     RECT  45.35 1.33 45.79 82.67 ;
     RECT  45.79 2.73 50.35 82.67 ;
     RECT  50.35 2.73 50.79 84.07 ;
     RECT  50.79 2.73 55.35 82.67 ;
     RECT  55.35 1.33 55.79 82.67 ;
     RECT  55.79 2.73 60.35 82.67 ;
     RECT  60.35 2.73 60.79 84.07 ;
     RECT  60.79 2.73 65.35 82.67 ;
     RECT  65.35 1.33 65.79 82.67 ;
     RECT  65.79 2.73 70.35 82.67 ;
     RECT  70.35 2.73 70.79 84.07 ;
     RECT  70.79 2.73 75.35 82.67 ;
     RECT  75.35 1.33 75.79 82.67 ;
     RECT  75.79 2.73 80.35 82.67 ;
     RECT  80.35 2.73 80.79 84.07 ;
    LAYER metal6 ;
     RECT  5.29 0 80.85 85 ;
  END
END enfasi
END LIBRARY
