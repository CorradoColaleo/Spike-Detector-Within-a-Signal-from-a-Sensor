`timescale 1ns/1ps
module top (input logic clk, rst,
            input logic enable, din,
            input logic signed [10:0] x,
            output logic spike);


endmodule

