VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

VIA via1_2_1120_340_1_3_300_300
  VIARULE Via1Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal1 via1 metal2 ;
  CUTSPACING 0.08 0.08 ;
  ENCLOSURE 0.035 0.05 0.035 0.035 ;
  ROWCOL 1 3 ;
END via1_2_1120_340_1_3_300_300

VIA via2_3_1120_340_1_3_320_320
  VIARULE Via2Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal2 via2 metal3 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.035 0.035 ;
  ROWCOL 1 3 ;
END via2_3_1120_340_1_3_320_320

VIA via3_4_1120_340_1_3_320_320
  VIARULE Via3Array-0 ;
  CUTSIZE 0.07 0.07 ;
  LAYERS metal3 via3 metal4 ;
  CUTSPACING 0.09 0.09 ;
  ENCLOSURE 0.035 0.035 0.035 0.035 ;
  ROWCOL 1 3 ;
END via3_4_1120_340_1_3_320_320

VIA via4_5_1120_340_1_2_600_600
  VIARULE Via4Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal4 via4 metal5 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0 0 ;
  ROWCOL 1 2 ;
END via4_5_1120_340_1_2_600_600

VIA via5_6_1120_340_1_2_600_600
  VIARULE Via5Array-0 ;
  CUTSIZE 0.14 0.14 ;
  LAYERS metal5 via5 metal6 ;
  CUTSPACING 0.16 0.16 ;
  ENCLOSURE 0 0 0.06 0 ;
  ROWCOL 1 2 ;
END via5_6_1120_340_1_2_600_600

MACRO iir
  FOREIGN iir 0 0 ;
  CLASS BLOCK ;
  SIZE 75 BY 75 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  59.72 74.93 59.79 75 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.875 0.07 21.945 ;
    END
  END rst
  PIN x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  16.4 74.93 16.47 75 ;
    END
  END x[0]
  PIN x[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  74.93 63.595 75 63.665 ;
    END
  END x[10]
  PIN x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  74.93 42.315 75 42.385 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  74.93 21.035 75 21.105 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  74.16 74.93 74.23 75 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  58.58 0 58.65 0.07 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 32.515 0.07 32.585 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 11.235 0.07 11.305 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  73.02 0 73.09 0.07 ;
    END
  END x[7]
  PIN x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  0.82 0 0.89 0.07 ;
    END
  END x[8]
  PIN x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  15.26 0 15.33 0.07 ;
    END
  END x[9]
  PIN z[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  30.84 74.93 30.91 75 ;
    END
  END z[0]
  PIN z[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  74.93 10.395 75 10.465 ;
    END
  END z[10]
  PIN z[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  29.7 0 29.77 0.07 ;
    END
  END z[1]
  PIN z[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  1.96 74.93 2.03 75 ;
    END
  END z[2]
  PIN z[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  74.93 52.955 75 53.025 ;
    END
  END z[3]
  PIN z[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 53.795 0.07 53.865 ;
    END
  END z[4]
  PIN z[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  45.28 74.93 45.35 75 ;
    END
  END z[5]
  PIN z[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT  44.14 0 44.21 0.07 ;
    END
  END z[6]
  PIN z[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 43.155 0.07 43.225 ;
    END
  END z[7]
  PIN z[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 64.435 0.07 64.505 ;
    END
  END z[8]
  PIN z[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  74.93 31.675 75 31.745 ;
    END
  END z[9]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal6 ;
        RECT  65.29 74.86 65.85 75 ;
        RECT  65.29 0 65.85 0.14 ;
        RECT  55.29 74.86 55.85 75 ;
        RECT  55.29 0 55.85 0.14 ;
        RECT  45.29 74.86 45.85 75 ;
        RECT  45.29 0 45.85 0.14 ;
        RECT  35.29 74.86 35.85 75 ;
        RECT  35.29 0 35.85 0.14 ;
        RECT  25.29 74.86 25.85 75 ;
        RECT  25.29 0 25.85 0.14 ;
        RECT  15.29 74.86 15.85 75 ;
        RECT  15.29 0 15.85 0.14 ;
        RECT  5.29 74.86 5.85 75 ;
        RECT  5.29 0 5.85 0.14 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal6 ;
        RECT  70.29 74.86 70.85 75 ;
        RECT  70.29 0 70.85 0.14 ;
        RECT  60.29 74.86 60.85 75 ;
        RECT  60.29 0 60.85 0.14 ;
        RECT  50.29 74.86 50.85 75 ;
        RECT  50.29 0 50.85 0.14 ;
        RECT  40.29 74.86 40.85 75 ;
        RECT  40.29 0 40.85 0.14 ;
        RECT  30.29 74.86 30.85 75 ;
        RECT  30.29 0 30.85 0.14 ;
        RECT  20.29 74.86 20.85 75 ;
        RECT  20.29 0 20.85 0.14 ;
        RECT  10.29 74.86 10.85 75 ;
        RECT  10.29 0 10.85 0.14 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
     RECT  0.57 1.315 0.82 74.285 ;
     RECT  0.82 0.035 1.96 74.285 ;
     RECT  1.96 0.035 16.21 74.725 ;
     RECT  16.21 0.035 26.54 74.865 ;
     RECT  26.54 0.035 32.17 74.585 ;
     RECT  32.17 0.035 32.81 74.865 ;
     RECT  32.81 0.175 34.9 74.865 ;
     RECT  34.9 0.875 37.18 74.865 ;
     RECT  37.18 0.875 37.75 74.585 ;
     RECT  37.75 0.875 38.32 74.445 ;
     RECT  38.32 1.315 41.1 74.445 ;
     RECT  41.1 1.315 43.19 74.585 ;
     RECT  43.19 1.315 43.38 74.725 ;
     RECT  43.38 1.315 44.14 74.865 ;
     RECT  44.14 0.035 58.08 74.865 ;
     RECT  58.08 0.875 62.45 74.865 ;
     RECT  62.45 1.315 73.66 74.865 ;
     RECT  73.66 1.315 74.48 74.285 ;
     RECT  74.48 46.935 74.8 47.005 ;
    LAYER metal2 ;
     RECT  29.89 0 31.29 0.035 ;
     RECT  29.7 0.035 32.81 0.175 ;
     RECT  0.82 0.035 0.89 0.245 ;
     RECT  29.7 0.175 34.9 0.875 ;
     RECT  58.01 0.035 58.65 0.875 ;
     RECT  56.87 0.875 62.45 1.015 ;
     RECT  15.26 0.035 15.33 1.155 ;
     RECT  21.15 0.875 24.83 1.155 ;
     RECT  56.68 1.015 62.45 1.155 ;
     RECT  13.74 1.155 24.83 1.33 ;
     RECT  44.14 0.035 44.21 1.33 ;
     RECT  50.98 1.155 62.45 1.33 ;
     RECT  5.34 1.33 5.8 1.715 ;
     RECT  29.7 0.875 38.32 1.715 ;
     RECT  50.98 1.33 65.8 1.715 ;
     RECT  5.34 1.715 9.25 1.855 ;
     RECT  13.74 1.33 25.8 1.855 ;
     RECT  29.7 1.715 39.84 1.855 ;
     RECT  44.14 1.33 45.8 1.855 ;
     RECT  5.34 1.855 25.8 1.995 ;
     RECT  29.7 1.855 45.8 1.995 ;
     RECT  50.98 1.715 68.91 1.995 ;
     RECT  73.02 0.035 73.09 1.995 ;
     RECT  5.34 1.995 73.09 2.555 ;
     RECT  5.34 2.555 73.28 3.605 ;
     RECT  5.34 3.605 72.71 6.615 ;
     RECT  4.81 6.615 72.71 7.595 ;
     RECT  4.81 7.595 73.47 7.735 ;
     RECT  4.24 7.735 73.47 8.715 ;
     RECT  3.67 8.715 73.47 9.135 ;
     RECT  3.67 9.135 74.42 10.395 ;
     RECT  3.67 10.395 74.99 11.935 ;
     RECT  2.53 11.935 74.99 15.995 ;
     RECT  2.34 15.995 74.99 17.115 ;
     RECT  1.58 17.115 74.99 18.375 ;
     RECT  0.63 18.375 74.99 21.945 ;
     RECT  0.82 21.945 74.99 24.185 ;
     RECT  1.01 24.185 74.99 32.375 ;
     RECT  0.82 32.375 74.99 32.445 ;
     RECT  1.39 32.445 74.99 39.655 ;
     RECT  1.2 39.655 74.99 40.075 ;
     RECT  1.01 40.075 74.99 40.845 ;
     RECT  1.58 40.845 74.99 45.255 ;
     RECT  1.01 45.255 74.99 45.745 ;
     RECT  1.77 45.745 74.99 46.865 ;
     RECT  2.34 46.865 74.99 47.005 ;
     RECT  2.34 47.005 73.85 51.135 ;
     RECT  2.15 51.135 73.85 51.275 ;
     RECT  1.39 51.275 73.85 51.975 ;
     RECT  1.2 51.975 73.85 52.045 ;
     RECT  1.58 52.045 73.85 52.465 ;
     RECT  1.77 52.465 73.85 55.125 ;
     RECT  1.96 55.125 73.85 56.245 ;
     RECT  2.34 56.245 73.85 56.805 ;
     RECT  2.72 56.805 73.85 58.065 ;
     RECT  2.91 58.065 73.85 58.555 ;
     RECT  2.91 58.555 74.23 60.865 ;
     RECT  4.24 60.865 74.23 61.005 ;
     RECT  5.34 61.005 74.23 66.115 ;
     RECT  4.81 66.115 74.23 67.935 ;
     RECT  3.67 67.935 74.23 68.845 ;
     RECT  4.43 68.845 74.23 69.545 ;
     RECT  5.34 69.545 74.23 73.745 ;
     RECT  5.34 73.745 31.1 74.27 ;
     RECT  35.34 73.745 74.23 74.27 ;
     RECT  6.9 74.27 31.1 74.445 ;
     RECT  36.16 74.27 63.21 74.445 ;
     RECT  67.13 74.27 74.23 74.445 ;
     RECT  6.9 74.445 6.97 74.585 ;
     RECT  11.46 74.445 18.94 74.585 ;
     RECT  36.16 74.445 45.35 74.585 ;
     RECT  69.98 74.445 74.23 74.585 ;
     RECT  12.6 74.585 16.47 74.725 ;
     RECT  26.09 74.445 31.1 74.725 ;
     RECT  43.19 74.585 45.35 74.725 ;
     RECT  16.21 74.725 16.47 74.865 ;
     RECT  29.89 74.725 31.1 74.865 ;
     RECT  37.11 74.585 37.18 74.865 ;
     RECT  43.38 74.725 45.35 74.865 ;
     RECT  50.41 74.445 62.26 74.865 ;
     RECT  71.69 74.585 74.23 74.865 ;
     RECT  1.96 74.655 2.03 74.965 ;
     RECT  16.4 74.865 16.47 74.965 ;
     RECT  29.89 74.865 30.91 74.965 ;
     RECT  45.28 74.865 45.35 74.965 ;
     RECT  59.72 74.865 59.79 74.965 ;
     RECT  74.16 74.865 74.23 74.965 ;
     RECT  29.89 74.965 30.72 75 ;
    LAYER metal3 ;
     RECT  0 11.375 0.035 12.005 ;
     RECT  0 22.015 0.035 22.645 ;
     RECT  0 43.295 0.035 43.645 ;
     RECT  0 64.155 0.035 64.365 ;
     RECT  0.035 11.235 0.13 12.005 ;
     RECT  0.035 64.155 0.13 64.505 ;
     RECT  0.035 43.155 1.01 43.645 ;
     RECT  0.035 32.515 1.2 32.585 ;
     RECT  1.01 38.255 1.2 38.325 ;
     RECT  1.01 43.155 1.2 45.325 ;
     RECT  1.2 42.875 1.39 45.465 ;
     RECT  1.39 18.655 1.58 18.725 ;
     RECT  0.035 21.875 1.58 22.645 ;
     RECT  1.39 27.475 1.58 27.545 ;
     RECT  1.2 32.515 1.58 32.865 ;
     RECT  1.58 27.055 1.77 27.545 ;
     RECT  1.58 32.515 1.77 33.145 ;
     RECT  1.2 38.255 1.77 38.745 ;
     RECT  1.39 42.455 1.77 45.465 ;
     RECT  0.035 53.795 1.77 53.865 ;
     RECT  1.77 27.055 1.96 34.405 ;
     RECT  1.96 25.935 2.15 34.405 ;
     RECT  1.77 38.255 2.15 46.865 ;
     RECT  2.15 25.935 2.34 46.865 ;
     RECT  2.15 50.855 2.34 50.925 ;
     RECT  1.77 53.795 2.34 54.705 ;
     RECT  0.13 11.935 2.53 12.005 ;
     RECT  2.34 25.935 2.53 55.265 ;
     RECT  2.53 25.935 2.72 56.805 ;
     RECT  1.58 17.115 2.91 18.725 ;
     RECT  1.58 21.875 2.91 23.065 ;
     RECT  2.72 25.935 3.1 56.945 ;
     RECT  3.67 8.715 3.86 8.785 ;
     RECT  2.53 11.935 4.05 13.545 ;
     RECT  2.91 17.115 4.05 23.065 ;
     RECT  3.86 8.715 4.24 9.065 ;
     RECT  3.67 68.775 4.43 68.845 ;
     RECT  4.05 11.935 4.62 23.065 ;
     RECT  3.1 25.935 4.62 61.005 ;
     RECT  4.24 7.735 4.81 9.065 ;
     RECT  4.62 11.935 4.81 61.005 ;
     RECT  0.13 64.155 4.81 64.225 ;
     RECT  4.43 68.775 4.81 69.545 ;
     RECT  4.81 6.615 5.34 61.005 ;
     RECT  4.81 64.155 5.34 69.545 ;
     RECT  5.34 1.33 5.8 74.27 ;
     RECT  5.8 1.995 8.87 73.885 ;
     RECT  8.87 1.995 10.39 73.745 ;
     RECT  10.39 1.995 10.465 73.605 ;
     RECT  10.465 1.855 10.77 73.605 ;
     RECT  10.77 1.855 10.8 72.87 ;
     RECT  10.8 1.855 13.93 72.205 ;
     RECT  13.93 1.855 15.34 73.605 ;
     RECT  15.34 1.33 15.8 74.27 ;
     RECT  15.8 2.135 21.53 73.605 ;
     RECT  21.53 1.995 24.19 73.605 ;
     RECT  24.19 1.995 25.34 73.885 ;
     RECT  25.34 1.33 25.8 74.27 ;
     RECT  25.8 1.995 27.11 74.025 ;
     RECT  27.11 1.995 30.08 73.885 ;
     RECT  30.08 1.855 31.03 73.885 ;
     RECT  31.03 1.855 32.24 74.865 ;
     RECT  32.24 1.855 35.34 73.325 ;
     RECT  35.34 1.33 35.8 74.27 ;
     RECT  35.8 1.855 36.73 74.27 ;
     RECT  36.73 1.855 41.93 74.445 ;
     RECT  41.93 2.135 45.34 74.445 ;
     RECT  45.34 1.33 45.8 74.445 ;
     RECT  45.8 8.855 46.11 74.445 ;
     RECT  45.8 1.995 48.7 4.725 ;
     RECT  46.11 8.855 48.7 73.605 ;
     RECT  48.7 1.995 48.96 73.605 ;
     RECT  48.96 2.275 50.03 73.605 ;
     RECT  50.03 2.275 53.71 74.865 ;
     RECT  53.71 2.275 54.21 74.725 ;
     RECT  54.21 2.135 55.34 74.725 ;
     RECT  55.34 1.33 55.8 74.725 ;
     RECT  55.8 1.995 55.99 74.725 ;
     RECT  55.99 1.995 59.53 70.945 ;
     RECT  59.53 1.995 59.72 71.085 ;
     RECT  55.99 74.515 59.72 74.725 ;
     RECT  59.72 1.995 60.36 74.725 ;
     RECT  60.36 2.135 63.52 74.725 ;
     RECT  63.52 1.995 63.97 74.725 ;
     RECT  63.97 1.995 65.34 74.27 ;
     RECT  65.34 1.33 65.8 74.27 ;
     RECT  65.8 1.995 68.53 52.185 ;
     RECT  65.8 55.195 69.79 72.345 ;
     RECT  68.53 2.135 70.34 52.185 ;
     RECT  69.79 55.195 70.34 73.605 ;
     RECT  70.34 2.135 70.8 73.605 ;
     RECT  70.8 60.795 70.81 73.605 ;
     RECT  70.81 67.795 71.19 73.605 ;
     RECT  70.8 2.135 71.38 35.665 ;
     RECT  71.38 5.775 71.76 35.665 ;
     RECT  71.38 2.135 71.88 2.625 ;
     RECT  70.81 60.795 71.95 64.785 ;
     RECT  70.8 38.955 72.33 45.605 ;
     RECT  71.95 60.795 72.33 63.665 ;
     RECT  71.76 5.775 72.52 35.525 ;
     RECT  71.19 67.795 72.52 73.465 ;
     RECT  72.52 6.335 72.71 21.105 ;
     RECT  72.33 39.935 72.71 45.605 ;
     RECT  72.52 67.795 72.71 72.205 ;
     RECT  72.71 17.815 72.9 21.105 ;
     RECT  72.71 39.935 72.9 44.205 ;
     RECT  72.71 67.795 72.9 68.005 ;
     RECT  71.88 1.995 73.09 2.625 ;
     RECT  72.52 23.975 73.09 35.525 ;
     RECT  72.9 41.195 73.09 44.205 ;
     RECT  72.33 63.035 73.09 63.665 ;
     RECT  72.71 70.875 73.09 72.205 ;
     RECT  73.09 2.555 73.28 2.625 ;
     RECT  72.9 18.655 73.28 21.105 ;
     RECT  73.09 70.875 73.28 72.065 ;
     RECT  72.71 6.335 73.47 14.945 ;
     RECT  73.09 29.575 73.47 35.525 ;
     RECT  73.28 70.875 73.47 70.945 ;
     RECT  73.28 20.335 73.66 21.105 ;
     RECT  73.09 23.975 73.66 26.005 ;
     RECT  73.47 29.575 73.66 33.145 ;
     RECT  70.8 51.975 73.66 53.585 ;
     RECT  72.9 67.795 73.66 67.865 ;
     RECT  73.47 9.135 73.85 14.945 ;
     RECT  73.66 31.675 73.85 33.145 ;
     RECT  73.66 24.255 74.04 26.005 ;
     RECT  73.85 31.675 74.04 33.005 ;
     RECT  73.66 20.895 74.05 21.105 ;
     RECT  73.85 14.875 74.23 14.945 ;
     RECT  74.04 25.935 74.23 26.005 ;
     RECT  73.85 9.135 74.42 10.465 ;
     RECT  73.09 42.315 74.8 44.205 ;
     RECT  74.42 10.395 74.965 10.465 ;
     RECT  74.05 21.035 74.965 21.105 ;
     RECT  74.04 31.675 74.965 31.745 ;
     RECT  74.8 42.315 74.965 42.385 ;
     RECT  73.66 51.975 74.965 53.025 ;
     RECT  73.09 63.595 74.965 63.665 ;
     RECT  74.965 51.975 75 52.885 ;
    LAYER metal4 ;
     RECT  35.34 1.33 35.8 1.96 ;
     RECT  5.34 1.33 5.8 2.73 ;
     RECT  15.34 1.33 15.8 2.73 ;
     RECT  25.34 1.33 25.8 2.73 ;
     RECT  35.025 1.96 35.8 2.73 ;
     RECT  45.34 1.33 45.8 2.73 ;
     RECT  55.34 1.33 55.8 2.73 ;
     RECT  65.34 1.33 65.8 2.73 ;
     RECT  5.34 2.73 70.8 16.94 ;
     RECT  4.785 16.94 70.8 25.62 ;
     RECT  5.34 25.62 70.8 32.06 ;
     RECT  5.34 32.06 72.685 35.7 ;
     RECT  4.785 35.7 72.685 35.98 ;
     RECT  4.225 35.98 72.685 36.68 ;
     RECT  3.945 36.68 72.685 40.04 ;
     RECT  3.945 40.04 70.8 44.66 ;
     RECT  2.545 44.66 70.8 49.7 ;
     RECT  4.785 49.7 70.8 55.58 ;
     RECT  5.34 55.58 70.8 72.87 ;
     RECT  5.34 72.87 5.8 74.27 ;
     RECT  15.34 72.87 15.8 74.27 ;
     RECT  25.34 72.87 25.8 74.27 ;
     RECT  35.34 72.87 35.8 74.27 ;
     RECT  45.34 72.87 45.8 74.27 ;
     RECT  55.34 72.87 55.8 74.27 ;
     RECT  63.865 72.87 65.8 74.27 ;
     RECT  63.865 74.27 64.005 74.76 ;
    LAYER metal5 ;
     RECT  5.35 1.33 5.79 74.27 ;
     RECT  5.79 2.73 15.35 72.87 ;
     RECT  15.35 1.33 15.79 74.27 ;
     RECT  15.79 2.73 25.35 72.87 ;
     RECT  25.35 1.33 25.79 74.27 ;
     RECT  25.79 2.73 35.35 72.87 ;
     RECT  35.35 1.33 35.79 74.27 ;
     RECT  35.79 2.73 45.35 72.87 ;
     RECT  45.35 1.33 45.79 74.27 ;
     RECT  45.79 2.73 55.35 72.87 ;
     RECT  55.35 1.33 55.79 74.27 ;
     RECT  55.79 2.73 65.35 72.87 ;
     RECT  65.35 1.33 65.79 74.27 ;
     RECT  65.79 2.73 70.79 72.87 ;
    LAYER metal6 ;
     RECT  5.29 0 70.85 75 ;
  END
END iir
END LIBRARY
