module top (clk,
    din,
    enable,
    rst,
    spike,
    x);
 input clk;
 input din;
 input enable;
 input rst;
 output spike;
 input [10:0] x;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire \blocco3.m1.soglia[0] ;
 wire \blocco3.m1.soglia[10] ;
 wire \blocco3.m1.soglia[11] ;
 wire \blocco3.m1.soglia[1] ;
 wire \blocco3.m1.soglia[2] ;
 wire \blocco3.m1.soglia[3] ;
 wire \blocco3.m1.soglia[4] ;
 wire \blocco3.m1.soglia[5] ;
 wire \blocco3.m1.soglia[6] ;
 wire \blocco3.m1.soglia[7] ;
 wire \blocco3.m1.soglia[8] ;
 wire \blocco3.m1.soglia[9] ;
 wire \blocco3.m2.q[0] ;
 wire \blocco3.m2.q[10] ;
 wire \blocco3.m2.q[11] ;
 wire \blocco3.m2.q[1] ;
 wire \blocco3.m2.q[2] ;
 wire \blocco3.m2.q[3] ;
 wire \blocco3.m2.q[4] ;
 wire \blocco3.m2.q[5] ;
 wire \blocco3.m2.q[6] ;
 wire \blocco3.m2.q[7] ;
 wire \blocco3.m2.q[8] ;
 wire \blocco3.m2.q[9] ;
 wire \blocco3.m2.stato_corrente[0] ;
 wire \blocco3.m2.stato_corrente[1] ;
 wire \blocco3.m2.stato_corrente[2] ;
 wire \output_iir[0] ;
 wire \output_iir[10] ;
 wire \output_iir[1] ;
 wire \output_iir[2] ;
 wire \output_iir[3] ;
 wire \output_iir[4] ;
 wire \output_iir[5] ;
 wire \output_iir[6] ;
 wire \output_iir[7] ;
 wire \output_iir[8] ;
 wire \output_iir[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire clk_regs;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_1_0__leaf_clk_regs;
 wire clknet_1_1__leaf_clk_regs;
 wire delaynet_0_my_clock;
 wire delaynet_1_my_clock;
 wire delaynet_2_my_clock;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;

 INV_X1 _110_ (.A(net9),
    .ZN(_045_));
 NAND2_X1 _111_ (.A1(net39),
    .A2(_045_),
    .ZN(_046_));
 NOR2_X1 _112_ (.A1(\blocco3.m2.stato_corrente[1] ),
    .A2(_046_),
    .ZN(spike));
 XOR2_X1 _113_ (.A(\blocco3.m1.soglia[11] ),
    .B(\blocco3.m2.q[11] ),
    .Z(_047_));
 XOR2_X1 _114_ (.A(\blocco3.m1.soglia[10] ),
    .B(\blocco3.m2.q[10] ),
    .Z(_048_));
 NOR2_X1 _115_ (.A1(_047_),
    .A2(_048_),
    .ZN(_049_));
 XOR2_X1 _116_ (.A(\blocco3.m1.soglia[9] ),
    .B(\blocco3.m2.q[9] ),
    .Z(_050_));
 XOR2_X1 _117_ (.A(\blocco3.m1.soglia[8] ),
    .B(\blocco3.m2.q[8] ),
    .Z(_051_));
 NOR2_X1 _118_ (.A1(_050_),
    .A2(_051_),
    .ZN(_052_));
 XOR2_X1 _119_ (.A(\blocco3.m1.soglia[7] ),
    .B(\blocco3.m2.q[7] ),
    .Z(_053_));
 XOR2_X1 _120_ (.A(\blocco3.m1.soglia[6] ),
    .B(\blocco3.m2.q[6] ),
    .Z(_054_));
 NOR2_X1 _121_ (.A1(_053_),
    .A2(_054_),
    .ZN(_055_));
 XOR2_X1 _122_ (.A(\blocco3.m1.soglia[5] ),
    .B(\blocco3.m2.q[5] ),
    .Z(_056_));
 XOR2_X1 _123_ (.A(\blocco3.m1.soglia[4] ),
    .B(\blocco3.m2.q[4] ),
    .Z(_057_));
 NOR2_X1 _124_ (.A1(_056_),
    .A2(_057_),
    .ZN(_058_));
 NAND4_X1 _125_ (.A1(_049_),
    .A2(_052_),
    .A3(_055_),
    .A4(_058_),
    .ZN(_059_));
 XOR2_X1 _126_ (.A(\blocco3.m1.soglia[3] ),
    .B(\blocco3.m2.q[3] ),
    .Z(_060_));
 XOR2_X1 _127_ (.A(\blocco3.m1.soglia[2] ),
    .B(\blocco3.m2.q[2] ),
    .Z(_061_));
 NOR2_X1 _128_ (.A1(_060_),
    .A2(_061_),
    .ZN(_062_));
 INV_X1 _129_ (.A(net12),
    .ZN(_063_));
 NOR2_X1 _130_ (.A1(_063_),
    .A2(\blocco3.m2.q[1] ),
    .ZN(_064_));
 XOR2_X1 _131_ (.A(\blocco3.m1.soglia[1] ),
    .B(\blocco3.m2.q[1] ),
    .Z(_065_));
 INV_X1 _132_ (.A(net21),
    .ZN(_066_));
 AOI21_X1 _133_ (.A(_065_),
    .B1(\blocco3.m2.q[0] ),
    .B2(_066_),
    .ZN(_067_));
 OAI21_X1 _134_ (.A(_062_),
    .B1(_064_),
    .B2(_067_),
    .ZN(_068_));
 INV_X1 _135_ (.A(net15),
    .ZN(_069_));
 NOR3_X1 _136_ (.A1(_069_),
    .A2(\blocco3.m2.q[2] ),
    .A3(_060_),
    .ZN(_070_));
 INV_X1 _137_ (.A(\blocco3.m2.q[3] ),
    .ZN(_071_));
 AOI21_X1 _138_ (.A(_070_),
    .B1(_071_),
    .B2(\blocco3.m1.soglia[3] ),
    .ZN(_072_));
 AOI21_X1 _139_ (.A(_059_),
    .B1(_068_),
    .B2(_072_),
    .ZN(_073_));
 INV_X1 _140_ (.A(net33),
    .ZN(_074_));
 NOR2_X1 _141_ (.A1(_074_),
    .A2(\blocco3.m2.q[9] ),
    .ZN(_075_));
 INV_X1 _142_ (.A(net36),
    .ZN(_076_));
 NOR3_X1 _143_ (.A1(_076_),
    .A2(\blocco3.m2.q[8] ),
    .A3(_050_),
    .ZN(_077_));
 OAI21_X1 _144_ (.A(_049_),
    .B1(_075_),
    .B2(_077_),
    .ZN(_078_));
 INV_X1 _145_ (.A(net18),
    .ZN(_079_));
 NOR3_X1 _146_ (.A1(_079_),
    .A2(\blocco3.m2.q[10] ),
    .A3(_047_),
    .ZN(_080_));
 INV_X1 _147_ (.A(net61),
    .ZN(_081_));
 AOI21_X1 _148_ (.A(_080_),
    .B1(_081_),
    .B2(\blocco3.m1.soglia[11] ),
    .ZN(_082_));
 NAND2_X1 _149_ (.A1(_078_),
    .A2(_082_),
    .ZN(_083_));
 NAND2_X1 _150_ (.A1(_049_),
    .A2(_052_),
    .ZN(_084_));
 INV_X1 _151_ (.A(net27),
    .ZN(_085_));
 NOR2_X1 _152_ (.A1(_085_),
    .A2(\blocco3.m2.q[5] ),
    .ZN(_086_));
 INV_X1 _153_ (.A(net24),
    .ZN(_087_));
 NOR3_X1 _154_ (.A1(_087_),
    .A2(\blocco3.m2.q[4] ),
    .A3(_056_),
    .ZN(_088_));
 OAI21_X1 _155_ (.A(_055_),
    .B1(_086_),
    .B2(_088_),
    .ZN(_089_));
 INV_X1 _156_ (.A(net30),
    .ZN(_090_));
 NOR3_X1 _157_ (.A1(_090_),
    .A2(\blocco3.m2.q[6] ),
    .A3(_053_),
    .ZN(_091_));
 INV_X1 _158_ (.A(\blocco3.m2.q[7] ),
    .ZN(_092_));
 AOI21_X1 _159_ (.A(_091_),
    .B1(_092_),
    .B2(\blocco3.m1.soglia[7] ),
    .ZN(_093_));
 AOI21_X1 _160_ (.A(_084_),
    .B1(_089_),
    .B2(_093_),
    .ZN(_094_));
 NOR4_X1 _161_ (.A1(_047_),
    .A2(_073_),
    .A3(_083_),
    .A4(_094_),
    .ZN(_095_));
 XOR2_X1 _162_ (.A(\blocco3.m1.soglia[0] ),
    .B(\blocco3.m2.q[0] ),
    .Z(_016_));
 NOR3_X1 _163_ (.A1(_059_),
    .A2(_065_),
    .A3(_016_),
    .ZN(_017_));
 AOI221_X1 _164_ (.A(_095_),
    .B1(_017_),
    .B2(_062_),
    .C1(_081_),
    .C2(\blocco3.m1.soglia[11] ),
    .ZN(_018_));
 OAI211_X1 _165_ (.A(net1),
    .B(net48),
    .C1(net9),
    .C2(_018_),
    .ZN(_019_));
 NOR2_X1 _166_ (.A1(net59),
    .A2(_045_),
    .ZN(_020_));
 OAI21_X1 _167_ (.A(_020_),
    .B1(net1),
    .B2(net39),
    .ZN(_021_));
 MUX2_X1 _168_ (.A(_046_),
    .B(_021_),
    .S(_018_),
    .Z(_022_));
 AOI21_X1 _169_ (.A(rst),
    .B1(net10),
    .B2(_022_),
    .ZN(_015_));
 NAND2_X1 _170_ (.A1(net1),
    .A2(_020_),
    .ZN(_023_));
 OR2_X1 _171_ (.A1(_018_),
    .A2(_023_),
    .ZN(_024_));
 AND3_X1 _172_ (.A1(net1),
    .A2(\blocco3.m2.stato_corrente[1] ),
    .A3(_045_),
    .ZN(_025_));
 AND2_X1 _173_ (.A1(net39),
    .A2(_020_),
    .ZN(_026_));
 AOI21_X1 _174_ (.A(_025_),
    .B1(_018_),
    .B2(net40),
    .ZN(_027_));
 AOI21_X1 _175_ (.A(rst),
    .B1(_024_),
    .B2(net41),
    .ZN(_014_));
 INV_X1 _176_ (.A(rst),
    .ZN(_028_));
 MUX2_X1 _177_ (.A(_045_),
    .B(_020_),
    .S(_018_),
    .Z(_029_));
 AND3_X1 _178_ (.A1(_028_),
    .A2(net47),
    .A3(_029_),
    .ZN(_013_));
 OAI21_X1 _179_ (.A(_028_),
    .B1(net33),
    .B2(enable),
    .ZN(_030_));
 AOI21_X1 _180_ (.A(_030_),
    .B1(enable),
    .B2(net37),
    .ZN(_012_));
 OAI21_X1 _181_ (.A(_028_),
    .B1(net36),
    .B2(enable),
    .ZN(_031_));
 INV_X1 _182_ (.A(net3),
    .ZN(_032_));
 AOI21_X1 _183_ (.A(_031_),
    .B1(net4),
    .B2(enable),
    .ZN(_011_));
 OAI21_X1 _184_ (.A(_028_),
    .B1(enable),
    .B2(net3),
    .ZN(_033_));
 AOI21_X1 _185_ (.A(_033_),
    .B1(net31),
    .B2(enable),
    .ZN(_010_));
 OAI21_X1 _186_ (.A(_028_),
    .B1(enable),
    .B2(net30),
    .ZN(_034_));
 AOI21_X1 _187_ (.A(_034_),
    .B1(net28),
    .B2(enable),
    .ZN(_009_));
 OAI21_X1 _188_ (.A(_028_),
    .B1(enable),
    .B2(net27),
    .ZN(_035_));
 AOI21_X1 _189_ (.A(_035_),
    .B1(net25),
    .B2(enable),
    .ZN(_008_));
 OAI21_X1 _190_ (.A(_028_),
    .B1(enable),
    .B2(net24),
    .ZN(_036_));
 INV_X1 _191_ (.A(net6),
    .ZN(_037_));
 AOI21_X1 _192_ (.A(_036_),
    .B1(net7),
    .B2(enable),
    .ZN(_007_));
 OAI21_X1 _193_ (.A(_028_),
    .B1(enable),
    .B2(net6),
    .ZN(_038_));
 AOI21_X1 _194_ (.A(_038_),
    .B1(net16),
    .B2(enable),
    .ZN(_006_));
 OAI21_X1 _195_ (.A(_028_),
    .B1(enable),
    .B2(net15),
    .ZN(_039_));
 AOI21_X1 _196_ (.A(_039_),
    .B1(net13),
    .B2(enable),
    .ZN(_005_));
 OAI21_X1 _197_ (.A(_028_),
    .B1(enable),
    .B2(net12),
    .ZN(_040_));
 AOI21_X1 _198_ (.A(_040_),
    .B1(net22),
    .B2(enable),
    .ZN(_004_));
 OAI21_X1 _199_ (.A(_028_),
    .B1(enable),
    .B2(net44),
    .ZN(_041_));
 AOI21_X1 _200_ (.A(net45),
    .B1(net19),
    .B2(enable),
    .ZN(_003_));
 OAI21_X1 _201_ (.A(_028_),
    .B1(enable),
    .B2(net18),
    .ZN(_042_));
 AOI21_X1 _202_ (.A(_042_),
    .B1(enable),
    .B2(net34),
    .ZN(_002_));
 OAI21_X1 _203_ (.A(_028_),
    .B1(enable),
    .B2(net21),
    .ZN(_043_));
 INV_X1 _204_ (.A(din),
    .ZN(_044_));
 AOI21_X1 _205_ (.A(_043_),
    .B1(_044_),
    .B2(enable),
    .ZN(_001_));
 iir blocco1 (.clk(clknet_1_0__leaf_clk),
    .rst(rst),
    .x({x[10],
    x[9],
    x[8],
    x[7],
    x[6],
    x[5],
    x[4],
    x[3],
    x[2],
    x[1],
    x[0]}),
    .z({\output_iir[10] ,
    \output_iir[9] ,
    \output_iir[8] ,
    \output_iir[7] ,
    \output_iir[6] ,
    \output_iir[5] ,
    \output_iir[4] ,
    \output_iir[3] ,
    \output_iir[2] ,
    \output_iir[1] ,
    \output_iir[0] }));
 enfasi blocco2 (.clk(clknet_1_1__leaf_clk),
    .rst(rst),
    .q({\blocco3.m2.q[11] ,
    \blocco3.m2.q[10] ,
    \blocco3.m2.q[9] ,
    \blocco3.m2.q[8] ,
    \blocco3.m2.q[7] ,
    \blocco3.m2.q[6] ,
    \blocco3.m2.q[5] ,
    \blocco3.m2.q[4] ,
    \blocco3.m2.q[3] ,
    \blocco3.m2.q[2] ,
    \blocco3.m2.q[1] ,
    \blocco3.m2.q[0] }),
    .z({\output_iir[10] ,
    \output_iir[9] ,
    \output_iir[8] ,
    \output_iir[7] ,
    \output_iir[6] ,
    \output_iir[5] ,
    \output_iir[4] ,
    \output_iir[3] ,
    \output_iir[2] ,
    \output_iir[1] ,
    \output_iir[0] }));
 DFF_X1 \blocco3.m1.soglia[0]$_SDFFE_PP0P_  (.D(_001_),
    .CK(clknet_1_1__leaf_clk_regs),
    .Q(\blocco3.m1.soglia[0] ),
    .QN(_109_));
 DFF_X1 \blocco3.m1.soglia[10]$_SDFFE_PP0P_  (.D(net35),
    .CK(clknet_1_0__leaf_clk_regs),
    .Q(\blocco3.m1.soglia[10] ),
    .QN(_108_));
 DFF_X1 \blocco3.m1.soglia[11]$_SDFFE_PP0P_  (.D(net20),
    .CK(clknet_1_0__leaf_clk_regs),
    .Q(\blocco3.m1.soglia[11] ),
    .QN(_107_));
 DFF_X1 \blocco3.m1.soglia[1]$_SDFFE_PP0P_  (.D(net23),
    .CK(clknet_1_1__leaf_clk_regs),
    .Q(\blocco3.m1.soglia[1] ),
    .QN(_106_));
 DFF_X1 \blocco3.m1.soglia[2]$_SDFFE_PP0P_  (.D(net14),
    .CK(clknet_1_1__leaf_clk_regs),
    .Q(\blocco3.m1.soglia[2] ),
    .QN(_105_));
 DFF_X1 \blocco3.m1.soglia[3]$_SDFFE_PP0P_  (.D(net17),
    .CK(clknet_1_1__leaf_clk_regs),
    .Q(\blocco3.m1.soglia[3] ),
    .QN(_104_));
 DFF_X1 \blocco3.m1.soglia[4]$_SDFFE_PP0P_  (.D(net8),
    .CK(clknet_1_1__leaf_clk_regs),
    .Q(\blocco3.m1.soglia[4] ),
    .QN(_103_));
 DFF_X1 \blocco3.m1.soglia[5]$_SDFFE_PP0P_  (.D(net26),
    .CK(clknet_1_1__leaf_clk_regs),
    .Q(\blocco3.m1.soglia[5] ),
    .QN(_102_));
 DFF_X1 \blocco3.m1.soglia[6]$_SDFFE_PP0P_  (.D(net29),
    .CK(clknet_1_0__leaf_clk_regs),
    .Q(\blocco3.m1.soglia[6] ),
    .QN(_101_));
 DFF_X1 \blocco3.m1.soglia[7]$_SDFFE_PP0P_  (.D(net32),
    .CK(clknet_1_0__leaf_clk_regs),
    .Q(\blocco3.m1.soglia[7] ),
    .QN(_100_));
 DFF_X1 \blocco3.m1.soglia[8]$_SDFFE_PP0P_  (.D(net5),
    .CK(clknet_1_0__leaf_clk_regs),
    .Q(\blocco3.m1.soglia[8] ),
    .QN(_099_));
 DFF_X1 \blocco3.m1.soglia[9]$_SDFFE_PP0P_  (.D(net38),
    .CK(clknet_1_0__leaf_clk_regs),
    .Q(\blocco3.m1.soglia[9] ),
    .QN(_098_));
 DFF_X1 \blocco3.m2.stato_corrente[0]$_SDFF_PP0_  (.D(net2),
    .CK(clknet_1_1__leaf_clk_regs),
    .Q(\blocco3.m2.stato_corrente[0] ),
    .QN(_097_));
 DFF_X1 \blocco3.m2.stato_corrente[1]$_SDFF_PP0_  (.D(net42),
    .CK(clknet_1_1__leaf_clk_regs),
    .Q(\blocco3.m2.stato_corrente[1] ),
    .QN(_096_));
 DFF_X1 \blocco3.m2.stato_corrente[2]$_SDFF_PP0_  (.D(net11),
    .CK(clknet_1_1__leaf_clk_regs),
    .Q(\blocco3.m2.stato_corrente[2] ),
    .QN(_000_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_2_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_2_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_2_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_2_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_3_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_3_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_3_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_3_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_3_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_3_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_3_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_3_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_3_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_3_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_3_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_3_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_3_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_3_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_3_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_3_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_3_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_3_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_3_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_3_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_3_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_3_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_3_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_3_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_3_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_3_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_3_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_3_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_3_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_3_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_3_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_3_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_3_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_3_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_3_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_3_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_3_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_3_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_3_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_3_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_3_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_3_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_3_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_3_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_3_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_3_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_3_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_3_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_3_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_3_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_3_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_3_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_3_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_3_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_3_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_3_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_3_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_1_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_1_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_1_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_1_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_1_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_1_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_1_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_1_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_1_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_1_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_1_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_1_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_1_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_1_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_1_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_1_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_1_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_1_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_1_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_1_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_1_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_1_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_1_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_1_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_1_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_1_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_1_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_1_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_1_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_1_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_1_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_1_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_1_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_1_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_1_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Left_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Left_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Left_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Left_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Left_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Left_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Left_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Left_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Left_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Left_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Left_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Left_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Left_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Left_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Left_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Left_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Left_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Left_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Left_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Left_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Left_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Left_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Left_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Left_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Left_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Left_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Left_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Left_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_1_Left_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_2_Left_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_2_Left_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_2_Left_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_2_Left_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_2_Left_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_2_Left_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_2_Left_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_2_Left_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_2_Left_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_2_Left_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_2_Left_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_2_Left_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_2_Left_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_2_Left_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_2_Left_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_2_Left_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_2_Left_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_2_Left_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_2_Left_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_2_Left_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_2_Left_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_2_Left_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_2_Left_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_2_Left_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_2_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_2_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_2_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_2_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_2_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_2_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_2_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_2_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_1_Right_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_1_Right_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_1_Right_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_1_Right_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_1_Right_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_1_Right_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_1_Right_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_1_Right_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_1_Right_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_1_Right_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_1_Right_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_1_Right_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_1_Right_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_1_Right_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_1_Right_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_1_Right_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_1_Right_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_1_Right_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_1_Right_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_1_Right_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_1_Right_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_1_Right_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_1_Right_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_1_Right_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_1_Right_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_1_Right_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_1_Right_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_1_Right_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_1_Right_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_1_Right_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_1_Right_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_1_Right_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Right_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Right_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Right_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Right_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Right_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Right_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Right_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Right_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Right_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Right_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Right_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Right_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Right_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Right_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Right_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Right_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Right_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Right_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Right_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Right_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Right_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Right_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Right_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Right_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Right_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_2_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_2_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_2_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_2_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_3_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_3_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_3_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_3_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_3_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_3_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_3_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_3_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_3_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_3_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_3_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_3_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_3_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_3_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_3_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_3_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_3_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_3_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_3_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_3_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_3_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_3_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_3_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_3_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_3_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_3_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_3_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_3_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_3_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_3_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_3_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_3_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_3_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_3_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_3_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_3_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_3_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_3_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_3_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_3_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_3_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_3_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_3_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_3_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_3_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_3_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_3_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_3_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_3_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_3_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_3_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_3_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_3_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_3_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_3_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_3_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_3_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_1_Right_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_1_Right_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_1_Right_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Right_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Right_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Right_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Right_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_1_Right_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_2_Right_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_2_Right_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_2_Right_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_2_Right_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_2_Right_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_2_Right_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_2_Right_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_2_Right_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_2_Right_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_2_Right_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_2_Right_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_2_Right_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_2_Right_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_2_Right_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_2_Right_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_2_Right_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_2_Right_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_2_Right_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_2_Right_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_2_Right_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_2_Right_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_2_Right_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_2_Right_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_2_Right_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_2_Right_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_2_Right_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_2_Right_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_2_Right_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_2_Right_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_2_Right_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_2_Right_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_2_Right_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Right_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Right_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Right_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Right_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Right_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Right_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Right_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Right_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Right_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Right_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Right_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Right_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Right_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Right_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Right_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Right_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Right_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Right_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Right_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Right_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Right_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Right_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Right_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Right_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Right_389 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_390 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_391 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_392 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_393 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_394 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_395 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_396 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_397 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_398 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_399 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_400 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_401 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_402 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_403 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_404 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_405 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_406 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_407 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_408 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_409 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_410 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_411 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_412 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_413 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_414 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_415 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_416 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_417 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_418 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_419 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_420 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_421 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_422 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_1_423 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_1_424 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_1_425 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_1_426 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_1_427 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_1_428 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_1_429 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_1_430 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_1_431 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_1_432 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_1_433 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_1_434 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_1_435 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_1_436 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_1_437 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_1_438 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_1_439 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_1_440 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_1_441 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_1_442 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_1_443 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_1_444 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_1_445 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_1_446 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_1_447 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_1_448 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_1_449 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_450 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_451 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_452 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_453 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_454 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_455 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_456 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_457 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_458 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_459 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_460 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_461 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_462 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_463 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_464 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_465 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_466 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_467 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_468 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_469 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_470 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_471 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_472 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_473 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_474 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_475 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_476 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_477 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_478 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_479 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_480 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_481 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_482 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_1_483 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_1_484 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_1_485 ();
 CLKBUF_X1 hold1 (.A(net46),
    .Z(net1));
 CLKBUF_X1 hold2 (.A(_013_),
    .Z(net2));
 CLKBUF_X1 hold3 (.A(net55),
    .Z(net3));
 CLKBUF_X1 hold4 (.A(_032_),
    .Z(net4));
 CLKBUF_X1 hold5 (.A(_011_),
    .Z(net5));
 CLKBUF_X1 hold6 (.A(net57),
    .Z(net6));
 CLKBUF_X1 hold7 (.A(_037_),
    .Z(net7));
 CLKBUF_X1 hold8 (.A(_007_),
    .Z(net8));
 CLKBUF_X1 hold9 (.A(\blocco3.m2.stato_corrente[0] ),
    .Z(net9));
 CLKBUF_X1 hold10 (.A(_019_),
    .Z(net10));
 CLKBUF_X1 hold11 (.A(net62),
    .Z(net11));
 CLKBUF_X1 hold12 (.A(net53),
    .Z(net12));
 CLKBUF_X1 hold13 (.A(_063_),
    .Z(net13));
 CLKBUF_X1 hold14 (.A(_005_),
    .Z(net14));
 CLKBUF_X1 hold15 (.A(net51),
    .Z(net15));
 CLKBUF_X1 hold16 (.A(_069_),
    .Z(net16));
 CLKBUF_X1 hold17 (.A(_006_),
    .Z(net17));
 CLKBUF_X1 hold18 (.A(net56),
    .Z(net18));
 CLKBUF_X1 hold19 (.A(_079_),
    .Z(net19));
 CLKBUF_X1 hold20 (.A(_003_),
    .Z(net20));
 CLKBUF_X1 hold21 (.A(net43),
    .Z(net21));
 CLKBUF_X1 hold22 (.A(_066_),
    .Z(net22));
 CLKBUF_X1 hold23 (.A(_004_),
    .Z(net23));
 CLKBUF_X1 hold24 (.A(net54),
    .Z(net24));
 CLKBUF_X1 hold25 (.A(_087_),
    .Z(net25));
 CLKBUF_X1 hold26 (.A(_008_),
    .Z(net26));
 CLKBUF_X1 hold27 (.A(net52),
    .Z(net27));
 CLKBUF_X1 hold28 (.A(_085_),
    .Z(net28));
 CLKBUF_X1 hold29 (.A(_009_),
    .Z(net29));
 CLKBUF_X1 hold30 (.A(net60),
    .Z(net30));
 CLKBUF_X1 hold31 (.A(_090_),
    .Z(net31));
 CLKBUF_X1 hold32 (.A(_010_),
    .Z(net32));
 CLKBUF_X1 hold33 (.A(net49),
    .Z(net33));
 CLKBUF_X1 hold34 (.A(_074_),
    .Z(net34));
 CLKBUF_X1 hold35 (.A(_002_),
    .Z(net35));
 CLKBUF_X1 hold36 (.A(net50),
    .Z(net36));
 CLKBUF_X1 hold37 (.A(_076_),
    .Z(net37));
 CLKBUF_X1 hold38 (.A(_012_),
    .Z(net38));
 CLKBUF_X1 hold39 (.A(\blocco3.m2.stato_corrente[2] ),
    .Z(net39));
 CLKBUF_X1 hold40 (.A(_026_),
    .Z(net40));
 CLKBUF_X1 hold41 (.A(_027_),
    .Z(net41));
 CLKBUF_X1 hold42 (.A(_014_),
    .Z(net42));
 CLKBUF_X1 hold43 (.A(net58),
    .Z(net43));
 CLKBUF_X1 hold44 (.A(\blocco3.m1.soglia[11] ),
    .Z(net44));
 CLKBUF_X1 hold45 (.A(_041_),
    .Z(net45));
 CLKBUF_X1 hold46 (.A(_000_),
    .Z(net46));
 CLKBUF_X1 hold47 (.A(net1),
    .Z(net47));
 CLKBUF_X1 hold48 (.A(\blocco3.m2.stato_corrente[1] ),
    .Z(net48));
 CLKBUF_X1 hold49 (.A(\blocco3.m1.soglia[9] ),
    .Z(net49));
 CLKBUF_X1 hold50 (.A(\blocco3.m1.soglia[8] ),
    .Z(net50));
 CLKBUF_X1 hold51 (.A(\blocco3.m1.soglia[2] ),
    .Z(net51));
 CLKBUF_X1 hold52 (.A(\blocco3.m1.soglia[5] ),
    .Z(net52));
 CLKBUF_X1 hold53 (.A(\blocco3.m1.soglia[1] ),
    .Z(net53));
 CLKBUF_X1 hold54 (.A(\blocco3.m1.soglia[4] ),
    .Z(net54));
 CLKBUF_X1 hold55 (.A(\blocco3.m1.soglia[7] ),
    .Z(net55));
 CLKBUF_X1 hold56 (.A(\blocco3.m1.soglia[10] ),
    .Z(net56));
 CLKBUF_X1 hold57 (.A(\blocco3.m1.soglia[3] ),
    .Z(net57));
 BUF_X8 clkbuf_regs_0_my_clock (.A(clk),
    .Z(delaynet_0_my_clock));
 BUF_X8 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 BUF_X8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 BUF_X8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 BUF_X1 clkload0 (.A(clknet_1_1__leaf_clk));
 BUF_X8 clkbuf_0_clk_regs (.A(clk_regs),
    .Z(clknet_0_clk_regs));
 BUF_X8 clkbuf_1_0__f_clk_regs (.A(clknet_0_clk_regs),
    .Z(clknet_1_0__leaf_clk_regs));
 BUF_X8 clkbuf_1_1__f_clk_regs (.A(clknet_0_clk_regs),
    .Z(clknet_1_1__leaf_clk_regs));
 INV_X2 clkload1 (.A(clknet_1_0__leaf_clk_regs));
 BUF_X8 delaybuf_0_my_clock (.A(delaynet_0_my_clock),
    .Z(delaynet_1_my_clock));
 BUF_X8 delaybuf_1_my_clock (.A(delaynet_1_my_clock),
    .Z(delaynet_2_my_clock));
 BUF_X8 delaybuf_2_my_clock (.A(delaynet_2_my_clock),
    .Z(clk_regs));
 CLKBUF_X1 hold58 (.A(\blocco3.m1.soglia[0] ),
    .Z(net58));
 CLKBUF_X1 hold59 (.A(\blocco3.m2.stato_corrente[1] ),
    .Z(net59));
 CLKBUF_X1 hold60 (.A(\blocco3.m1.soglia[6] ),
    .Z(net60));
 CLKBUF_X1 hold61 (.A(\blocco3.m2.q[11] ),
    .Z(net61));
 CLKBUF_X1 hold62 (.A(_015_),
    .Z(net62));
 FILLCELL_X32 FILLER_0_0_1 ();
 FILLCELL_X32 FILLER_0_0_33 ();
 FILLCELL_X16 FILLER_0_0_65 ();
 FILLCELL_X8 FILLER_0_0_81 ();
 FILLCELL_X32 FILLER_0_0_90 ();
 FILLCELL_X32 FILLER_0_0_122 ();
 FILLCELL_X16 FILLER_0_0_154 ();
 FILLCELL_X8 FILLER_0_0_170 ();
 FILLCELL_X32 FILLER_0_0_179 ();
 FILLCELL_X32 FILLER_0_0_211 ();
 FILLCELL_X16 FILLER_0_0_243 ();
 FILLCELL_X8 FILLER_0_0_259 ();
 FILLCELL_X32 FILLER_0_0_268 ();
 FILLCELL_X32 FILLER_0_0_300 ();
 FILLCELL_X16 FILLER_0_0_332 ();
 FILLCELL_X8 FILLER_0_0_348 ();
 FILLCELL_X32 FILLER_0_0_357 ();
 FILLCELL_X32 FILLER_0_0_389 ();
 FILLCELL_X16 FILLER_0_0_421 ();
 FILLCELL_X8 FILLER_0_0_437 ();
 FILLCELL_X32 FILLER_0_0_446 ();
 FILLCELL_X32 FILLER_0_0_478 ();
 FILLCELL_X16 FILLER_0_0_510 ();
 FILLCELL_X8 FILLER_0_0_526 ();
 FILLCELL_X32 FILLER_0_0_535 ();
 FILLCELL_X32 FILLER_0_0_567 ();
 FILLCELL_X16 FILLER_0_0_599 ();
 FILLCELL_X8 FILLER_0_0_615 ();
 FILLCELL_X32 FILLER_0_0_624 ();
 FILLCELL_X32 FILLER_0_0_656 ();
 FILLCELL_X16 FILLER_0_0_688 ();
 FILLCELL_X8 FILLER_0_0_704 ();
 FILLCELL_X32 FILLER_0_0_713 ();
 FILLCELL_X32 FILLER_0_0_745 ();
 FILLCELL_X16 FILLER_0_0_777 ();
 FILLCELL_X8 FILLER_0_0_793 ();
 FILLCELL_X32 FILLER_0_0_802 ();
 FILLCELL_X32 FILLER_0_0_834 ();
 FILLCELL_X16 FILLER_0_0_866 ();
 FILLCELL_X8 FILLER_0_0_882 ();
 FILLCELL_X32 FILLER_0_0_891 ();
 FILLCELL_X32 FILLER_0_0_923 ();
 FILLCELL_X16 FILLER_0_0_955 ();
 FILLCELL_X8 FILLER_0_0_971 ();
 FILLCELL_X32 FILLER_0_0_980 ();
 FILLCELL_X32 FILLER_0_0_1012 ();
 FILLCELL_X2 FILLER_0_0_1044 ();
 FILLCELL_X32 FILLER_0_1_1 ();
 FILLCELL_X32 FILLER_0_1_33 ();
 FILLCELL_X32 FILLER_0_1_65 ();
 FILLCELL_X32 FILLER_0_1_97 ();
 FILLCELL_X32 FILLER_0_1_129 ();
 FILLCELL_X16 FILLER_0_1_161 ();
 FILLCELL_X1 FILLER_0_1_177 ();
 FILLCELL_X32 FILLER_0_1_179 ();
 FILLCELL_X32 FILLER_0_1_211 ();
 FILLCELL_X32 FILLER_0_1_243 ();
 FILLCELL_X32 FILLER_0_1_275 ();
 FILLCELL_X32 FILLER_0_1_307 ();
 FILLCELL_X16 FILLER_0_1_339 ();
 FILLCELL_X1 FILLER_0_1_355 ();
 FILLCELL_X32 FILLER_0_1_357 ();
 FILLCELL_X32 FILLER_0_1_389 ();
 FILLCELL_X32 FILLER_0_1_421 ();
 FILLCELL_X32 FILLER_0_1_453 ();
 FILLCELL_X32 FILLER_0_1_485 ();
 FILLCELL_X16 FILLER_0_1_517 ();
 FILLCELL_X1 FILLER_0_1_533 ();
 FILLCELL_X32 FILLER_0_1_535 ();
 FILLCELL_X32 FILLER_0_1_567 ();
 FILLCELL_X32 FILLER_0_1_599 ();
 FILLCELL_X32 FILLER_0_1_631 ();
 FILLCELL_X32 FILLER_0_1_663 ();
 FILLCELL_X16 FILLER_0_1_695 ();
 FILLCELL_X1 FILLER_0_1_711 ();
 FILLCELL_X32 FILLER_0_1_713 ();
 FILLCELL_X32 FILLER_0_1_745 ();
 FILLCELL_X32 FILLER_0_1_777 ();
 FILLCELL_X32 FILLER_0_1_809 ();
 FILLCELL_X32 FILLER_0_1_841 ();
 FILLCELL_X16 FILLER_0_1_873 ();
 FILLCELL_X1 FILLER_0_1_889 ();
 FILLCELL_X32 FILLER_0_1_891 ();
 FILLCELL_X32 FILLER_0_1_923 ();
 FILLCELL_X32 FILLER_0_1_955 ();
 FILLCELL_X32 FILLER_0_1_987 ();
 FILLCELL_X16 FILLER_0_1_1019 ();
 FILLCELL_X8 FILLER_0_1_1035 ();
 FILLCELL_X2 FILLER_0_1_1043 ();
 FILLCELL_X1 FILLER_0_1_1045 ();
 FILLCELL_X32 FILLER_0_2_1 ();
 FILLCELL_X32 FILLER_0_2_33 ();
 FILLCELL_X16 FILLER_0_2_65 ();
 FILLCELL_X8 FILLER_0_2_81 ();
 FILLCELL_X32 FILLER_0_2_90 ();
 FILLCELL_X32 FILLER_0_2_122 ();
 FILLCELL_X32 FILLER_0_2_154 ();
 FILLCELL_X32 FILLER_0_2_186 ();
 FILLCELL_X32 FILLER_0_2_218 ();
 FILLCELL_X16 FILLER_0_2_250 ();
 FILLCELL_X1 FILLER_0_2_266 ();
 FILLCELL_X32 FILLER_0_2_268 ();
 FILLCELL_X32 FILLER_0_2_300 ();
 FILLCELL_X32 FILLER_0_2_332 ();
 FILLCELL_X32 FILLER_0_2_364 ();
 FILLCELL_X32 FILLER_0_2_396 ();
 FILLCELL_X16 FILLER_0_2_428 ();
 FILLCELL_X1 FILLER_0_2_444 ();
 FILLCELL_X32 FILLER_0_2_446 ();
 FILLCELL_X32 FILLER_0_2_478 ();
 FILLCELL_X32 FILLER_0_2_510 ();
 FILLCELL_X32 FILLER_0_2_542 ();
 FILLCELL_X32 FILLER_0_2_574 ();
 FILLCELL_X16 FILLER_0_2_606 ();
 FILLCELL_X1 FILLER_0_2_622 ();
 FILLCELL_X32 FILLER_0_2_624 ();
 FILLCELL_X32 FILLER_0_2_656 ();
 FILLCELL_X32 FILLER_0_2_688 ();
 FILLCELL_X32 FILLER_0_2_720 ();
 FILLCELL_X32 FILLER_0_2_752 ();
 FILLCELL_X16 FILLER_0_2_784 ();
 FILLCELL_X1 FILLER_0_2_800 ();
 FILLCELL_X32 FILLER_0_2_802 ();
 FILLCELL_X32 FILLER_0_2_834 ();
 FILLCELL_X32 FILLER_0_2_866 ();
 FILLCELL_X32 FILLER_0_2_898 ();
 FILLCELL_X32 FILLER_0_2_930 ();
 FILLCELL_X16 FILLER_0_2_962 ();
 FILLCELL_X1 FILLER_0_2_978 ();
 FILLCELL_X32 FILLER_0_2_980 ();
 FILLCELL_X32 FILLER_0_2_1012 ();
 FILLCELL_X2 FILLER_0_2_1044 ();
 FILLCELL_X32 FILLER_0_3_1 ();
 FILLCELL_X32 FILLER_0_3_33 ();
 FILLCELL_X16 FILLER_0_3_65 ();
 FILLCELL_X8 FILLER_0_3_81 ();
 FILLCELL_X32 FILLER_0_3_90 ();
 FILLCELL_X32 FILLER_0_3_122 ();
 FILLCELL_X16 FILLER_0_3_154 ();
 FILLCELL_X8 FILLER_0_3_170 ();
 FILLCELL_X32 FILLER_0_3_179 ();
 FILLCELL_X32 FILLER_0_3_211 ();
 FILLCELL_X16 FILLER_0_3_243 ();
 FILLCELL_X8 FILLER_0_3_259 ();
 FILLCELL_X32 FILLER_0_3_268 ();
 FILLCELL_X32 FILLER_0_3_300 ();
 FILLCELL_X16 FILLER_0_3_332 ();
 FILLCELL_X8 FILLER_0_3_348 ();
 FILLCELL_X32 FILLER_0_3_357 ();
 FILLCELL_X32 FILLER_0_3_389 ();
 FILLCELL_X16 FILLER_0_3_421 ();
 FILLCELL_X8 FILLER_0_3_437 ();
 FILLCELL_X32 FILLER_0_3_446 ();
 FILLCELL_X32 FILLER_0_3_478 ();
 FILLCELL_X16 FILLER_0_3_510 ();
 FILLCELL_X8 FILLER_0_3_526 ();
 FILLCELL_X32 FILLER_0_3_535 ();
 FILLCELL_X32 FILLER_0_3_567 ();
 FILLCELL_X16 FILLER_0_3_599 ();
 FILLCELL_X8 FILLER_0_3_615 ();
 FILLCELL_X32 FILLER_0_3_624 ();
 FILLCELL_X32 FILLER_0_3_656 ();
 FILLCELL_X16 FILLER_0_3_688 ();
 FILLCELL_X8 FILLER_0_3_704 ();
 FILLCELL_X32 FILLER_0_3_713 ();
 FILLCELL_X8 FILLER_0_3_745 ();
 FILLCELL_X32 FILLER_0_3_756 ();
 FILLCELL_X8 FILLER_0_3_788 ();
 FILLCELL_X4 FILLER_0_3_796 ();
 FILLCELL_X1 FILLER_0_3_800 ();
 FILLCELL_X32 FILLER_0_3_802 ();
 FILLCELL_X32 FILLER_0_3_834 ();
 FILLCELL_X16 FILLER_0_3_866 ();
 FILLCELL_X8 FILLER_0_3_882 ();
 FILLCELL_X32 FILLER_0_3_891 ();
 FILLCELL_X32 FILLER_0_3_923 ();
 FILLCELL_X16 FILLER_0_3_955 ();
 FILLCELL_X8 FILLER_0_3_971 ();
 FILLCELL_X32 FILLER_0_3_980 ();
 FILLCELL_X32 FILLER_0_3_1012 ();
 FILLCELL_X2 FILLER_0_3_1044 ();
 FILLCELL_X32 FILLER_0_4_1 ();
 FILLCELL_X32 FILLER_0_4_33 ();
 FILLCELL_X16 FILLER_0_4_65 ();
 FILLCELL_X8 FILLER_0_4_81 ();
 FILLCELL_X32 FILLER_0_4_90 ();
 FILLCELL_X32 FILLER_0_4_122 ();
 FILLCELL_X32 FILLER_0_4_154 ();
 FILLCELL_X32 FILLER_0_4_186 ();
 FILLCELL_X32 FILLER_0_4_218 ();
 FILLCELL_X16 FILLER_0_4_250 ();
 FILLCELL_X1 FILLER_0_4_266 ();
 FILLCELL_X32 FILLER_0_4_268 ();
 FILLCELL_X32 FILLER_0_4_300 ();
 FILLCELL_X32 FILLER_0_4_332 ();
 FILLCELL_X32 FILLER_0_4_364 ();
 FILLCELL_X32 FILLER_0_4_396 ();
 FILLCELL_X16 FILLER_0_4_428 ();
 FILLCELL_X1 FILLER_0_4_444 ();
 FILLCELL_X32 FILLER_0_4_446 ();
 FILLCELL_X32 FILLER_0_4_478 ();
 FILLCELL_X16 FILLER_0_4_510 ();
 FILLCELL_X8 FILLER_0_4_526 ();
 FILLCELL_X2 FILLER_0_4_534 ();
 FILLCELL_X1 FILLER_0_4_536 ();
 FILLCELL_X32 FILLER_0_4_1008 ();
 FILLCELL_X4 FILLER_0_4_1040 ();
 FILLCELL_X2 FILLER_0_4_1044 ();
 FILLCELL_X32 FILLER_0_5_1 ();
 FILLCELL_X32 FILLER_0_5_33 ();
 FILLCELL_X32 FILLER_0_5_65 ();
 FILLCELL_X32 FILLER_0_5_97 ();
 FILLCELL_X32 FILLER_0_5_129 ();
 FILLCELL_X16 FILLER_0_5_161 ();
 FILLCELL_X1 FILLER_0_5_177 ();
 FILLCELL_X32 FILLER_0_5_179 ();
 FILLCELL_X32 FILLER_0_5_211 ();
 FILLCELL_X32 FILLER_0_5_243 ();
 FILLCELL_X32 FILLER_0_5_275 ();
 FILLCELL_X32 FILLER_0_5_307 ();
 FILLCELL_X16 FILLER_0_5_339 ();
 FILLCELL_X1 FILLER_0_5_355 ();
 FILLCELL_X32 FILLER_0_5_357 ();
 FILLCELL_X32 FILLER_0_5_389 ();
 FILLCELL_X32 FILLER_0_5_421 ();
 FILLCELL_X32 FILLER_0_5_453 ();
 FILLCELL_X32 FILLER_0_5_485 ();
 FILLCELL_X16 FILLER_0_5_517 ();
 FILLCELL_X1 FILLER_0_5_533 ();
 FILLCELL_X2 FILLER_0_5_535 ();
 FILLCELL_X32 FILLER_0_5_1008 ();
 FILLCELL_X4 FILLER_0_5_1040 ();
 FILLCELL_X2 FILLER_0_5_1044 ();
 FILLCELL_X32 FILLER_0_6_1 ();
 FILLCELL_X32 FILLER_0_6_33 ();
 FILLCELL_X16 FILLER_0_6_65 ();
 FILLCELL_X8 FILLER_0_6_81 ();
 FILLCELL_X32 FILLER_0_6_90 ();
 FILLCELL_X32 FILLER_0_6_122 ();
 FILLCELL_X32 FILLER_0_6_154 ();
 FILLCELL_X32 FILLER_0_6_186 ();
 FILLCELL_X32 FILLER_0_6_218 ();
 FILLCELL_X16 FILLER_0_6_250 ();
 FILLCELL_X1 FILLER_0_6_266 ();
 FILLCELL_X8 FILLER_0_6_268 ();
 FILLCELL_X4 FILLER_0_6_276 ();
 FILLCELL_X2 FILLER_0_6_280 ();
 FILLCELL_X1 FILLER_0_6_282 ();
 FILLCELL_X32 FILLER_0_6_296 ();
 FILLCELL_X32 FILLER_0_6_328 ();
 FILLCELL_X32 FILLER_0_6_360 ();
 FILLCELL_X32 FILLER_0_6_392 ();
 FILLCELL_X16 FILLER_0_6_424 ();
 FILLCELL_X4 FILLER_0_6_440 ();
 FILLCELL_X1 FILLER_0_6_444 ();
 FILLCELL_X32 FILLER_0_6_446 ();
 FILLCELL_X32 FILLER_0_6_478 ();
 FILLCELL_X16 FILLER_0_6_510 ();
 FILLCELL_X8 FILLER_0_6_526 ();
 FILLCELL_X2 FILLER_0_6_534 ();
 FILLCELL_X1 FILLER_0_6_536 ();
 FILLCELL_X32 FILLER_0_6_1008 ();
 FILLCELL_X4 FILLER_0_6_1040 ();
 FILLCELL_X2 FILLER_0_6_1044 ();
 FILLCELL_X32 FILLER_0_7_1 ();
 FILLCELL_X32 FILLER_0_7_33 ();
 FILLCELL_X16 FILLER_0_7_65 ();
 FILLCELL_X8 FILLER_0_7_81 ();
 FILLCELL_X32 FILLER_0_7_90 ();
 FILLCELL_X32 FILLER_0_7_122 ();
 FILLCELL_X16 FILLER_0_7_154 ();
 FILLCELL_X8 FILLER_0_7_170 ();
 FILLCELL_X32 FILLER_0_7_179 ();
 FILLCELL_X32 FILLER_0_7_211 ();
 FILLCELL_X16 FILLER_0_7_243 ();
 FILLCELL_X8 FILLER_0_7_259 ();
 FILLCELL_X32 FILLER_0_7_268 ();
 FILLCELL_X32 FILLER_0_7_300 ();
 FILLCELL_X16 FILLER_0_7_332 ();
 FILLCELL_X8 FILLER_0_7_348 ();
 FILLCELL_X32 FILLER_0_7_357 ();
 FILLCELL_X32 FILLER_0_7_389 ();
 FILLCELL_X16 FILLER_0_7_421 ();
 FILLCELL_X8 FILLER_0_7_437 ();
 FILLCELL_X32 FILLER_0_7_446 ();
 FILLCELL_X32 FILLER_0_7_478 ();
 FILLCELL_X16 FILLER_0_7_510 ();
 FILLCELL_X8 FILLER_0_7_526 ();
 FILLCELL_X2 FILLER_0_7_535 ();
 FILLCELL_X32 FILLER_0_7_1008 ();
 FILLCELL_X4 FILLER_0_7_1040 ();
 FILLCELL_X2 FILLER_0_7_1044 ();
 FILLCELL_X32 FILLER_0_8_1 ();
 FILLCELL_X4 FILLER_0_8_33 ();
 FILLCELL_X32 FILLER_0_8_456 ();
 FILLCELL_X32 FILLER_0_8_488 ();
 FILLCELL_X16 FILLER_0_8_520 ();
 FILLCELL_X1 FILLER_0_8_536 ();
 FILLCELL_X32 FILLER_0_8_1008 ();
 FILLCELL_X4 FILLER_0_8_1040 ();
 FILLCELL_X2 FILLER_0_8_1044 ();
 FILLCELL_X32 FILLER_0_9_1 ();
 FILLCELL_X4 FILLER_0_9_33 ();
 FILLCELL_X32 FILLER_0_9_456 ();
 FILLCELL_X32 FILLER_0_9_488 ();
 FILLCELL_X16 FILLER_0_9_520 ();
 FILLCELL_X1 FILLER_0_9_536 ();
 FILLCELL_X32 FILLER_0_9_1008 ();
 FILLCELL_X4 FILLER_0_9_1040 ();
 FILLCELL_X2 FILLER_0_9_1044 ();
 FILLCELL_X32 FILLER_0_10_1 ();
 FILLCELL_X4 FILLER_0_10_33 ();
 FILLCELL_X32 FILLER_0_10_456 ();
 FILLCELL_X32 FILLER_0_10_488 ();
 FILLCELL_X16 FILLER_0_10_520 ();
 FILLCELL_X1 FILLER_0_10_536 ();
 FILLCELL_X32 FILLER_0_10_1008 ();
 FILLCELL_X4 FILLER_0_10_1040 ();
 FILLCELL_X2 FILLER_0_10_1044 ();
 FILLCELL_X32 FILLER_0_11_1 ();
 FILLCELL_X4 FILLER_0_11_33 ();
 FILLCELL_X32 FILLER_0_11_456 ();
 FILLCELL_X32 FILLER_0_11_488 ();
 FILLCELL_X16 FILLER_0_11_520 ();
 FILLCELL_X1 FILLER_0_11_536 ();
 FILLCELL_X32 FILLER_0_11_1008 ();
 FILLCELL_X4 FILLER_0_11_1040 ();
 FILLCELL_X2 FILLER_0_11_1044 ();
 FILLCELL_X32 FILLER_0_12_1 ();
 FILLCELL_X4 FILLER_0_12_33 ();
 FILLCELL_X32 FILLER_0_12_456 ();
 FILLCELL_X32 FILLER_0_12_488 ();
 FILLCELL_X16 FILLER_0_12_520 ();
 FILLCELL_X1 FILLER_0_12_536 ();
 FILLCELL_X32 FILLER_0_12_1008 ();
 FILLCELL_X4 FILLER_0_12_1040 ();
 FILLCELL_X2 FILLER_0_12_1044 ();
 FILLCELL_X32 FILLER_0_13_1 ();
 FILLCELL_X4 FILLER_0_13_33 ();
 FILLCELL_X32 FILLER_0_13_456 ();
 FILLCELL_X32 FILLER_0_13_488 ();
 FILLCELL_X16 FILLER_0_13_520 ();
 FILLCELL_X1 FILLER_0_13_536 ();
 FILLCELL_X32 FILLER_0_13_1008 ();
 FILLCELL_X4 FILLER_0_13_1040 ();
 FILLCELL_X2 FILLER_0_13_1044 ();
 FILLCELL_X32 FILLER_0_14_1 ();
 FILLCELL_X4 FILLER_0_14_33 ();
 FILLCELL_X32 FILLER_0_14_456 ();
 FILLCELL_X32 FILLER_0_14_488 ();
 FILLCELL_X16 FILLER_0_14_520 ();
 FILLCELL_X1 FILLER_0_14_536 ();
 FILLCELL_X32 FILLER_0_14_1008 ();
 FILLCELL_X4 FILLER_0_14_1040 ();
 FILLCELL_X2 FILLER_0_14_1044 ();
 FILLCELL_X32 FILLER_0_15_1 ();
 FILLCELL_X4 FILLER_0_15_33 ();
 FILLCELL_X32 FILLER_0_15_456 ();
 FILLCELL_X32 FILLER_0_15_488 ();
 FILLCELL_X16 FILLER_0_15_520 ();
 FILLCELL_X1 FILLER_0_15_536 ();
 FILLCELL_X32 FILLER_0_15_1008 ();
 FILLCELL_X4 FILLER_0_15_1040 ();
 FILLCELL_X2 FILLER_0_15_1044 ();
 FILLCELL_X32 FILLER_0_16_1 ();
 FILLCELL_X4 FILLER_0_16_33 ();
 FILLCELL_X32 FILLER_0_16_456 ();
 FILLCELL_X32 FILLER_0_16_488 ();
 FILLCELL_X16 FILLER_0_16_520 ();
 FILLCELL_X1 FILLER_0_16_536 ();
 FILLCELL_X32 FILLER_0_16_1008 ();
 FILLCELL_X4 FILLER_0_16_1040 ();
 FILLCELL_X2 FILLER_0_16_1044 ();
 FILLCELL_X32 FILLER_0_17_1 ();
 FILLCELL_X4 FILLER_0_17_33 ();
 FILLCELL_X32 FILLER_0_17_456 ();
 FILLCELL_X32 FILLER_0_17_488 ();
 FILLCELL_X16 FILLER_0_17_520 ();
 FILLCELL_X1 FILLER_0_17_536 ();
 FILLCELL_X32 FILLER_0_17_1008 ();
 FILLCELL_X4 FILLER_0_17_1040 ();
 FILLCELL_X2 FILLER_0_17_1044 ();
 FILLCELL_X32 FILLER_0_18_1 ();
 FILLCELL_X4 FILLER_0_18_33 ();
 FILLCELL_X32 FILLER_0_18_456 ();
 FILLCELL_X32 FILLER_0_18_488 ();
 FILLCELL_X16 FILLER_0_18_520 ();
 FILLCELL_X1 FILLER_0_18_536 ();
 FILLCELL_X32 FILLER_0_18_1008 ();
 FILLCELL_X4 FILLER_0_18_1040 ();
 FILLCELL_X2 FILLER_0_18_1044 ();
 FILLCELL_X32 FILLER_0_19_1 ();
 FILLCELL_X4 FILLER_0_19_33 ();
 FILLCELL_X32 FILLER_0_19_456 ();
 FILLCELL_X32 FILLER_0_19_488 ();
 FILLCELL_X16 FILLER_0_19_520 ();
 FILLCELL_X1 FILLER_0_19_536 ();
 FILLCELL_X32 FILLER_0_19_1008 ();
 FILLCELL_X4 FILLER_0_19_1040 ();
 FILLCELL_X2 FILLER_0_19_1044 ();
 FILLCELL_X32 FILLER_0_20_1 ();
 FILLCELL_X4 FILLER_0_20_33 ();
 FILLCELL_X32 FILLER_0_20_456 ();
 FILLCELL_X32 FILLER_0_20_488 ();
 FILLCELL_X16 FILLER_0_20_520 ();
 FILLCELL_X1 FILLER_0_20_536 ();
 FILLCELL_X32 FILLER_0_20_1008 ();
 FILLCELL_X4 FILLER_0_20_1040 ();
 FILLCELL_X2 FILLER_0_20_1044 ();
 FILLCELL_X32 FILLER_0_21_1 ();
 FILLCELL_X4 FILLER_0_21_33 ();
 FILLCELL_X32 FILLER_0_21_456 ();
 FILLCELL_X32 FILLER_0_21_488 ();
 FILLCELL_X16 FILLER_0_21_520 ();
 FILLCELL_X1 FILLER_0_21_536 ();
 FILLCELL_X32 FILLER_0_21_1008 ();
 FILLCELL_X4 FILLER_0_21_1040 ();
 FILLCELL_X2 FILLER_0_21_1044 ();
 FILLCELL_X32 FILLER_0_22_1 ();
 FILLCELL_X4 FILLER_0_22_33 ();
 FILLCELL_X8 FILLER_0_22_456 ();
 FILLCELL_X1 FILLER_0_22_464 ();
 FILLCELL_X32 FILLER_0_22_478 ();
 FILLCELL_X16 FILLER_0_22_510 ();
 FILLCELL_X8 FILLER_0_22_526 ();
 FILLCELL_X2 FILLER_0_22_534 ();
 FILLCELL_X1 FILLER_0_22_536 ();
 FILLCELL_X32 FILLER_0_22_1008 ();
 FILLCELL_X4 FILLER_0_22_1040 ();
 FILLCELL_X2 FILLER_0_22_1044 ();
 FILLCELL_X32 FILLER_0_23_1 ();
 FILLCELL_X4 FILLER_0_23_33 ();
 FILLCELL_X16 FILLER_0_23_456 ();
 FILLCELL_X4 FILLER_0_23_472 ();
 FILLCELL_X32 FILLER_0_23_489 ();
 FILLCELL_X16 FILLER_0_23_521 ();
 FILLCELL_X32 FILLER_0_23_1008 ();
 FILLCELL_X4 FILLER_0_23_1040 ();
 FILLCELL_X2 FILLER_0_23_1044 ();
 FILLCELL_X32 FILLER_0_24_1 ();
 FILLCELL_X4 FILLER_0_24_33 ();
 FILLCELL_X16 FILLER_0_24_456 ();
 FILLCELL_X8 FILLER_0_24_472 ();
 FILLCELL_X2 FILLER_0_24_480 ();
 FILLCELL_X16 FILLER_0_24_495 ();
 FILLCELL_X8 FILLER_0_24_511 ();
 FILLCELL_X8 FILLER_0_24_527 ();
 FILLCELL_X2 FILLER_0_24_535 ();
 FILLCELL_X32 FILLER_0_24_1008 ();
 FILLCELL_X4 FILLER_0_24_1040 ();
 FILLCELL_X2 FILLER_0_24_1044 ();
 FILLCELL_X32 FILLER_0_25_1 ();
 FILLCELL_X4 FILLER_0_25_33 ();
 FILLCELL_X32 FILLER_0_25_456 ();
 FILLCELL_X16 FILLER_0_25_488 ();
 FILLCELL_X8 FILLER_0_25_504 ();
 FILLCELL_X2 FILLER_0_25_512 ();
 FILLCELL_X1 FILLER_0_25_520 ();
 FILLCELL_X8 FILLER_0_25_527 ();
 FILLCELL_X2 FILLER_0_25_535 ();
 FILLCELL_X32 FILLER_0_25_1008 ();
 FILLCELL_X4 FILLER_0_25_1040 ();
 FILLCELL_X2 FILLER_0_25_1044 ();
 FILLCELL_X32 FILLER_0_26_1 ();
 FILLCELL_X4 FILLER_0_26_33 ();
 FILLCELL_X32 FILLER_0_26_456 ();
 FILLCELL_X16 FILLER_0_26_488 ();
 FILLCELL_X4 FILLER_0_26_504 ();
 FILLCELL_X2 FILLER_0_26_508 ();
 FILLCELL_X1 FILLER_0_26_510 ();
 FILLCELL_X1 FILLER_0_26_520 ();
 FILLCELL_X8 FILLER_0_26_528 ();
 FILLCELL_X1 FILLER_0_26_536 ();
 FILLCELL_X32 FILLER_0_26_1008 ();
 FILLCELL_X4 FILLER_0_26_1040 ();
 FILLCELL_X2 FILLER_0_26_1044 ();
 FILLCELL_X32 FILLER_0_27_1 ();
 FILLCELL_X4 FILLER_0_27_33 ();
 FILLCELL_X32 FILLER_0_27_456 ();
 FILLCELL_X4 FILLER_0_27_488 ();
 FILLCELL_X2 FILLER_0_27_492 ();
 FILLCELL_X1 FILLER_0_27_494 ();
 FILLCELL_X1 FILLER_0_27_524 ();
 FILLCELL_X4 FILLER_0_27_531 ();
 FILLCELL_X2 FILLER_0_27_535 ();
 FILLCELL_X32 FILLER_0_27_1008 ();
 FILLCELL_X4 FILLER_0_27_1040 ();
 FILLCELL_X2 FILLER_0_27_1044 ();
 FILLCELL_X32 FILLER_0_28_1 ();
 FILLCELL_X4 FILLER_0_28_33 ();
 FILLCELL_X32 FILLER_0_28_456 ();
 FILLCELL_X4 FILLER_0_28_488 ();
 FILLCELL_X1 FILLER_0_28_525 ();
 FILLCELL_X4 FILLER_0_28_531 ();
 FILLCELL_X2 FILLER_0_28_535 ();
 FILLCELL_X32 FILLER_0_28_1008 ();
 FILLCELL_X4 FILLER_0_28_1040 ();
 FILLCELL_X2 FILLER_0_28_1044 ();
 FILLCELL_X32 FILLER_0_29_1 ();
 FILLCELL_X4 FILLER_0_29_33 ();
 FILLCELL_X32 FILLER_0_29_456 ();
 FILLCELL_X16 FILLER_0_29_488 ();
 FILLCELL_X4 FILLER_0_29_530 ();
 FILLCELL_X2 FILLER_0_29_534 ();
 FILLCELL_X1 FILLER_0_29_536 ();
 FILLCELL_X32 FILLER_0_29_1008 ();
 FILLCELL_X4 FILLER_0_29_1040 ();
 FILLCELL_X2 FILLER_0_29_1044 ();
 FILLCELL_X32 FILLER_0_30_1 ();
 FILLCELL_X4 FILLER_0_30_33 ();
 FILLCELL_X32 FILLER_0_30_456 ();
 FILLCELL_X8 FILLER_0_30_488 ();
 FILLCELL_X4 FILLER_0_30_496 ();
 FILLCELL_X2 FILLER_0_30_500 ();
 FILLCELL_X1 FILLER_0_30_502 ();
 FILLCELL_X1 FILLER_0_30_523 ();
 FILLCELL_X4 FILLER_0_30_530 ();
 FILLCELL_X2 FILLER_0_30_534 ();
 FILLCELL_X1 FILLER_0_30_536 ();
 FILLCELL_X32 FILLER_0_30_1008 ();
 FILLCELL_X4 FILLER_0_30_1040 ();
 FILLCELL_X2 FILLER_0_30_1044 ();
 FILLCELL_X32 FILLER_0_31_1 ();
 FILLCELL_X4 FILLER_0_31_33 ();
 FILLCELL_X32 FILLER_0_31_456 ();
 FILLCELL_X8 FILLER_0_31_488 ();
 FILLCELL_X4 FILLER_0_31_496 ();
 FILLCELL_X2 FILLER_0_31_528 ();
 FILLCELL_X4 FILLER_0_31_533 ();
 FILLCELL_X32 FILLER_0_31_1008 ();
 FILLCELL_X4 FILLER_0_31_1040 ();
 FILLCELL_X2 FILLER_0_31_1044 ();
 FILLCELL_X32 FILLER_0_32_1 ();
 FILLCELL_X4 FILLER_0_32_33 ();
 FILLCELL_X32 FILLER_0_32_456 ();
 FILLCELL_X8 FILLER_0_32_488 ();
 FILLCELL_X4 FILLER_0_32_496 ();
 FILLCELL_X2 FILLER_0_32_500 ();
 FILLCELL_X4 FILLER_0_32_521 ();
 FILLCELL_X1 FILLER_0_32_525 ();
 FILLCELL_X4 FILLER_0_32_530 ();
 FILLCELL_X2 FILLER_0_32_534 ();
 FILLCELL_X1 FILLER_0_32_536 ();
 FILLCELL_X32 FILLER_0_32_1008 ();
 FILLCELL_X4 FILLER_0_32_1040 ();
 FILLCELL_X2 FILLER_0_32_1044 ();
 FILLCELL_X32 FILLER_0_33_1 ();
 FILLCELL_X4 FILLER_0_33_33 ();
 FILLCELL_X32 FILLER_0_33_456 ();
 FILLCELL_X8 FILLER_0_33_488 ();
 FILLCELL_X4 FILLER_0_33_496 ();
 FILLCELL_X2 FILLER_0_33_500 ();
 FILLCELL_X1 FILLER_0_33_502 ();
 FILLCELL_X8 FILLER_0_33_516 ();
 FILLCELL_X4 FILLER_0_33_531 ();
 FILLCELL_X2 FILLER_0_33_535 ();
 FILLCELL_X32 FILLER_0_33_1008 ();
 FILLCELL_X4 FILLER_0_33_1040 ();
 FILLCELL_X2 FILLER_0_33_1044 ();
 FILLCELL_X32 FILLER_0_34_1 ();
 FILLCELL_X4 FILLER_0_34_33 ();
 FILLCELL_X32 FILLER_0_34_456 ();
 FILLCELL_X8 FILLER_0_34_488 ();
 FILLCELL_X2 FILLER_0_34_496 ();
 FILLCELL_X2 FILLER_0_34_522 ();
 FILLCELL_X1 FILLER_0_34_524 ();
 FILLCELL_X8 FILLER_0_34_528 ();
 FILLCELL_X1 FILLER_0_34_536 ();
 FILLCELL_X32 FILLER_0_34_1008 ();
 FILLCELL_X4 FILLER_0_34_1040 ();
 FILLCELL_X2 FILLER_0_34_1044 ();
 FILLCELL_X32 FILLER_0_35_1 ();
 FILLCELL_X4 FILLER_0_35_33 ();
 FILLCELL_X32 FILLER_0_35_456 ();
 FILLCELL_X4 FILLER_0_35_488 ();
 FILLCELL_X2 FILLER_0_35_492 ();
 FILLCELL_X1 FILLER_0_35_494 ();
 FILLCELL_X4 FILLER_0_35_497 ();
 FILLCELL_X1 FILLER_0_35_501 ();
 FILLCELL_X4 FILLER_0_35_533 ();
 FILLCELL_X32 FILLER_0_35_1008 ();
 FILLCELL_X4 FILLER_0_35_1040 ();
 FILLCELL_X2 FILLER_0_35_1044 ();
 FILLCELL_X32 FILLER_0_36_1 ();
 FILLCELL_X4 FILLER_0_36_33 ();
 FILLCELL_X16 FILLER_0_36_456 ();
 FILLCELL_X8 FILLER_0_36_472 ();
 FILLCELL_X2 FILLER_0_36_480 ();
 FILLCELL_X4 FILLER_0_36_485 ();
 FILLCELL_X1 FILLER_0_36_489 ();
 FILLCELL_X8 FILLER_0_36_494 ();
 FILLCELL_X4 FILLER_0_36_533 ();
 FILLCELL_X32 FILLER_0_36_1008 ();
 FILLCELL_X4 FILLER_0_36_1040 ();
 FILLCELL_X2 FILLER_0_36_1044 ();
 FILLCELL_X32 FILLER_0_37_1 ();
 FILLCELL_X4 FILLER_0_37_33 ();
 FILLCELL_X8 FILLER_0_37_456 ();
 FILLCELL_X4 FILLER_0_37_464 ();
 FILLCELL_X2 FILLER_0_37_468 ();
 FILLCELL_X1 FILLER_0_37_487 ();
 FILLCELL_X4 FILLER_0_37_505 ();
 FILLCELL_X2 FILLER_0_37_512 ();
 FILLCELL_X1 FILLER_0_37_514 ();
 FILLCELL_X2 FILLER_0_37_525 ();
 FILLCELL_X4 FILLER_0_37_532 ();
 FILLCELL_X1 FILLER_0_37_536 ();
 FILLCELL_X32 FILLER_0_37_1008 ();
 FILLCELL_X4 FILLER_0_37_1040 ();
 FILLCELL_X2 FILLER_0_37_1044 ();
 FILLCELL_X32 FILLER_0_38_1 ();
 FILLCELL_X4 FILLER_0_38_33 ();
 FILLCELL_X16 FILLER_0_38_456 ();
 FILLCELL_X8 FILLER_0_38_472 ();
 FILLCELL_X2 FILLER_0_38_500 ();
 FILLCELL_X1 FILLER_0_38_502 ();
 FILLCELL_X4 FILLER_0_38_533 ();
 FILLCELL_X32 FILLER_0_38_1008 ();
 FILLCELL_X4 FILLER_0_38_1040 ();
 FILLCELL_X2 FILLER_0_38_1044 ();
 FILLCELL_X32 FILLER_0_39_1 ();
 FILLCELL_X4 FILLER_0_39_33 ();
 FILLCELL_X8 FILLER_0_39_456 ();
 FILLCELL_X4 FILLER_0_39_464 ();
 FILLCELL_X2 FILLER_0_39_468 ();
 FILLCELL_X1 FILLER_0_39_506 ();
 FILLCELL_X4 FILLER_0_39_511 ();
 FILLCELL_X4 FILLER_0_39_532 ();
 FILLCELL_X1 FILLER_0_39_536 ();
 FILLCELL_X32 FILLER_0_39_1008 ();
 FILLCELL_X4 FILLER_0_39_1040 ();
 FILLCELL_X2 FILLER_0_39_1044 ();
 FILLCELL_X32 FILLER_0_40_1 ();
 FILLCELL_X4 FILLER_0_40_33 ();
 FILLCELL_X16 FILLER_0_40_456 ();
 FILLCELL_X2 FILLER_0_40_472 ();
 FILLCELL_X1 FILLER_0_40_510 ();
 FILLCELL_X1 FILLER_0_40_515 ();
 FILLCELL_X1 FILLER_0_40_522 ();
 FILLCELL_X4 FILLER_0_40_532 ();
 FILLCELL_X1 FILLER_0_40_536 ();
 FILLCELL_X32 FILLER_0_40_1008 ();
 FILLCELL_X4 FILLER_0_40_1040 ();
 FILLCELL_X2 FILLER_0_40_1044 ();
 FILLCELL_X32 FILLER_0_41_1 ();
 FILLCELL_X4 FILLER_0_41_33 ();
 FILLCELL_X16 FILLER_0_41_456 ();
 FILLCELL_X2 FILLER_0_41_472 ();
 FILLCELL_X2 FILLER_0_41_491 ();
 FILLCELL_X1 FILLER_0_41_493 ();
 FILLCELL_X2 FILLER_0_41_497 ();
 FILLCELL_X1 FILLER_0_41_499 ();
 FILLCELL_X1 FILLER_0_41_523 ();
 FILLCELL_X4 FILLER_0_41_530 ();
 FILLCELL_X2 FILLER_0_41_534 ();
 FILLCELL_X1 FILLER_0_41_536 ();
 FILLCELL_X32 FILLER_0_41_1008 ();
 FILLCELL_X4 FILLER_0_41_1040 ();
 FILLCELL_X2 FILLER_0_41_1044 ();
 FILLCELL_X32 FILLER_0_42_1 ();
 FILLCELL_X4 FILLER_0_42_33 ();
 FILLCELL_X16 FILLER_0_42_456 ();
 FILLCELL_X4 FILLER_0_42_472 ();
 FILLCELL_X2 FILLER_0_42_476 ();
 FILLCELL_X2 FILLER_0_42_485 ();
 FILLCELL_X1 FILLER_0_42_487 ();
 FILLCELL_X1 FILLER_0_42_491 ();
 FILLCELL_X4 FILLER_0_42_495 ();
 FILLCELL_X2 FILLER_0_42_499 ();
 FILLCELL_X8 FILLER_0_42_528 ();
 FILLCELL_X1 FILLER_0_42_536 ();
 FILLCELL_X32 FILLER_0_42_1008 ();
 FILLCELL_X4 FILLER_0_42_1040 ();
 FILLCELL_X2 FILLER_0_42_1044 ();
 FILLCELL_X32 FILLER_0_43_1 ();
 FILLCELL_X4 FILLER_0_43_33 ();
 FILLCELL_X16 FILLER_0_43_456 ();
 FILLCELL_X8 FILLER_0_43_472 ();
 FILLCELL_X4 FILLER_0_43_480 ();
 FILLCELL_X2 FILLER_0_43_484 ();
 FILLCELL_X1 FILLER_0_43_486 ();
 FILLCELL_X2 FILLER_0_43_514 ();
 FILLCELL_X2 FILLER_0_43_528 ();
 FILLCELL_X1 FILLER_0_43_530 ();
 FILLCELL_X2 FILLER_0_43_534 ();
 FILLCELL_X1 FILLER_0_43_536 ();
 FILLCELL_X32 FILLER_0_43_1008 ();
 FILLCELL_X4 FILLER_0_43_1040 ();
 FILLCELL_X2 FILLER_0_43_1044 ();
 FILLCELL_X32 FILLER_0_44_1 ();
 FILLCELL_X4 FILLER_0_44_33 ();
 FILLCELL_X16 FILLER_0_44_456 ();
 FILLCELL_X8 FILLER_0_44_472 ();
 FILLCELL_X4 FILLER_0_44_480 ();
 FILLCELL_X2 FILLER_0_44_488 ();
 FILLCELL_X2 FILLER_0_44_528 ();
 FILLCELL_X4 FILLER_0_44_532 ();
 FILLCELL_X1 FILLER_0_44_536 ();
 FILLCELL_X32 FILLER_0_44_1008 ();
 FILLCELL_X4 FILLER_0_44_1040 ();
 FILLCELL_X2 FILLER_0_44_1044 ();
 FILLCELL_X32 FILLER_0_45_1 ();
 FILLCELL_X4 FILLER_0_45_33 ();
 FILLCELL_X16 FILLER_0_45_456 ();
 FILLCELL_X8 FILLER_0_45_472 ();
 FILLCELL_X2 FILLER_0_45_480 ();
 FILLCELL_X1 FILLER_0_45_482 ();
 FILLCELL_X8 FILLER_0_45_489 ();
 FILLCELL_X4 FILLER_0_45_497 ();
 FILLCELL_X2 FILLER_0_45_508 ();
 FILLCELL_X1 FILLER_0_45_510 ();
 FILLCELL_X8 FILLER_0_45_529 ();
 FILLCELL_X32 FILLER_0_45_1008 ();
 FILLCELL_X4 FILLER_0_45_1040 ();
 FILLCELL_X2 FILLER_0_45_1044 ();
 FILLCELL_X32 FILLER_0_46_1 ();
 FILLCELL_X4 FILLER_0_46_33 ();
 FILLCELL_X16 FILLER_0_46_456 ();
 FILLCELL_X4 FILLER_0_46_472 ();
 FILLCELL_X2 FILLER_0_46_476 ();
 FILLCELL_X1 FILLER_0_46_478 ();
 FILLCELL_X8 FILLER_0_46_486 ();
 FILLCELL_X4 FILLER_0_46_494 ();
 FILLCELL_X8 FILLER_0_46_528 ();
 FILLCELL_X1 FILLER_0_46_536 ();
 FILLCELL_X32 FILLER_0_46_1008 ();
 FILLCELL_X4 FILLER_0_46_1040 ();
 FILLCELL_X2 FILLER_0_46_1044 ();
 FILLCELL_X32 FILLER_0_47_1 ();
 FILLCELL_X4 FILLER_0_47_33 ();
 FILLCELL_X16 FILLER_0_47_456 ();
 FILLCELL_X1 FILLER_0_47_472 ();
 FILLCELL_X1 FILLER_0_47_528 ();
 FILLCELL_X2 FILLER_0_47_535 ();
 FILLCELL_X32 FILLER_0_47_1008 ();
 FILLCELL_X4 FILLER_0_47_1040 ();
 FILLCELL_X2 FILLER_0_47_1044 ();
 FILLCELL_X32 FILLER_0_48_1 ();
 FILLCELL_X4 FILLER_0_48_33 ();
 FILLCELL_X32 FILLER_0_48_456 ();
 FILLCELL_X32 FILLER_0_48_488 ();
 FILLCELL_X16 FILLER_0_48_520 ();
 FILLCELL_X1 FILLER_0_48_536 ();
 FILLCELL_X32 FILLER_0_48_1008 ();
 FILLCELL_X4 FILLER_0_48_1040 ();
 FILLCELL_X2 FILLER_0_48_1044 ();
 FILLCELL_X32 FILLER_0_49_1 ();
 FILLCELL_X4 FILLER_0_49_33 ();
 FILLCELL_X32 FILLER_0_49_456 ();
 FILLCELL_X32 FILLER_0_49_488 ();
 FILLCELL_X16 FILLER_0_49_520 ();
 FILLCELL_X1 FILLER_0_49_536 ();
 FILLCELL_X32 FILLER_0_49_1008 ();
 FILLCELL_X4 FILLER_0_49_1040 ();
 FILLCELL_X2 FILLER_0_49_1044 ();
 FILLCELL_X32 FILLER_0_50_1 ();
 FILLCELL_X4 FILLER_0_50_33 ();
 FILLCELL_X32 FILLER_0_50_456 ();
 FILLCELL_X32 FILLER_0_50_488 ();
 FILLCELL_X16 FILLER_0_50_520 ();
 FILLCELL_X1 FILLER_0_50_536 ();
 FILLCELL_X32 FILLER_0_50_1008 ();
 FILLCELL_X4 FILLER_0_50_1040 ();
 FILLCELL_X2 FILLER_0_50_1044 ();
 FILLCELL_X32 FILLER_0_51_1 ();
 FILLCELL_X4 FILLER_0_51_33 ();
 FILLCELL_X32 FILLER_0_51_456 ();
 FILLCELL_X32 FILLER_0_51_488 ();
 FILLCELL_X4 FILLER_0_51_520 ();
 FILLCELL_X32 FILLER_0_51_1008 ();
 FILLCELL_X4 FILLER_0_51_1040 ();
 FILLCELL_X2 FILLER_0_51_1044 ();
 FILLCELL_X32 FILLER_0_52_1 ();
 FILLCELL_X4 FILLER_0_52_33 ();
 FILLCELL_X32 FILLER_0_52_456 ();
 FILLCELL_X32 FILLER_0_52_488 ();
 FILLCELL_X16 FILLER_0_52_520 ();
 FILLCELL_X1 FILLER_0_52_536 ();
 FILLCELL_X32 FILLER_0_52_1008 ();
 FILLCELL_X4 FILLER_0_52_1040 ();
 FILLCELL_X2 FILLER_0_52_1044 ();
 FILLCELL_X32 FILLER_0_53_1 ();
 FILLCELL_X4 FILLER_0_53_33 ();
 FILLCELL_X32 FILLER_0_53_456 ();
 FILLCELL_X32 FILLER_0_53_488 ();
 FILLCELL_X16 FILLER_0_53_520 ();
 FILLCELL_X1 FILLER_0_53_536 ();
 FILLCELL_X32 FILLER_0_53_1008 ();
 FILLCELL_X4 FILLER_0_53_1040 ();
 FILLCELL_X2 FILLER_0_53_1044 ();
 FILLCELL_X32 FILLER_0_54_1 ();
 FILLCELL_X4 FILLER_0_54_33 ();
 FILLCELL_X32 FILLER_0_54_456 ();
 FILLCELL_X32 FILLER_0_54_488 ();
 FILLCELL_X16 FILLER_0_54_520 ();
 FILLCELL_X1 FILLER_0_54_536 ();
 FILLCELL_X32 FILLER_0_54_1008 ();
 FILLCELL_X4 FILLER_0_54_1040 ();
 FILLCELL_X2 FILLER_0_54_1044 ();
 FILLCELL_X32 FILLER_0_55_1 ();
 FILLCELL_X4 FILLER_0_55_33 ();
 FILLCELL_X32 FILLER_0_55_456 ();
 FILLCELL_X32 FILLER_0_55_488 ();
 FILLCELL_X16 FILLER_0_55_520 ();
 FILLCELL_X1 FILLER_0_55_536 ();
 FILLCELL_X32 FILLER_0_55_1008 ();
 FILLCELL_X4 FILLER_0_55_1040 ();
 FILLCELL_X2 FILLER_0_55_1044 ();
 FILLCELL_X32 FILLER_0_56_1 ();
 FILLCELL_X4 FILLER_0_56_33 ();
 FILLCELL_X32 FILLER_0_56_456 ();
 FILLCELL_X32 FILLER_0_56_488 ();
 FILLCELL_X16 FILLER_0_56_520 ();
 FILLCELL_X1 FILLER_0_56_536 ();
 FILLCELL_X32 FILLER_0_56_1008 ();
 FILLCELL_X4 FILLER_0_56_1040 ();
 FILLCELL_X2 FILLER_0_56_1044 ();
 FILLCELL_X32 FILLER_0_57_1 ();
 FILLCELL_X4 FILLER_0_57_33 ();
 FILLCELL_X32 FILLER_0_57_456 ();
 FILLCELL_X32 FILLER_0_57_488 ();
 FILLCELL_X16 FILLER_0_57_520 ();
 FILLCELL_X1 FILLER_0_57_536 ();
 FILLCELL_X32 FILLER_0_57_1008 ();
 FILLCELL_X4 FILLER_0_57_1040 ();
 FILLCELL_X2 FILLER_0_57_1044 ();
 FILLCELL_X32 FILLER_0_58_1 ();
 FILLCELL_X4 FILLER_0_58_33 ();
 FILLCELL_X32 FILLER_0_58_456 ();
 FILLCELL_X32 FILLER_0_58_488 ();
 FILLCELL_X16 FILLER_0_58_520 ();
 FILLCELL_X1 FILLER_0_58_536 ();
 FILLCELL_X32 FILLER_0_58_1008 ();
 FILLCELL_X4 FILLER_0_58_1040 ();
 FILLCELL_X2 FILLER_0_58_1044 ();
 FILLCELL_X32 FILLER_0_59_1 ();
 FILLCELL_X4 FILLER_0_59_33 ();
 FILLCELL_X32 FILLER_0_59_456 ();
 FILLCELL_X32 FILLER_0_59_488 ();
 FILLCELL_X16 FILLER_0_59_520 ();
 FILLCELL_X1 FILLER_0_59_536 ();
 FILLCELL_X32 FILLER_0_59_1008 ();
 FILLCELL_X4 FILLER_0_59_1040 ();
 FILLCELL_X2 FILLER_0_59_1044 ();
 FILLCELL_X32 FILLER_0_60_1 ();
 FILLCELL_X4 FILLER_0_60_33 ();
 FILLCELL_X32 FILLER_0_60_456 ();
 FILLCELL_X32 FILLER_0_60_488 ();
 FILLCELL_X16 FILLER_0_60_520 ();
 FILLCELL_X1 FILLER_0_60_536 ();
 FILLCELL_X32 FILLER_0_60_1008 ();
 FILLCELL_X4 FILLER_0_60_1040 ();
 FILLCELL_X2 FILLER_0_60_1044 ();
 FILLCELL_X32 FILLER_0_61_1 ();
 FILLCELL_X4 FILLER_0_61_33 ();
 FILLCELL_X32 FILLER_0_61_456 ();
 FILLCELL_X32 FILLER_0_61_488 ();
 FILLCELL_X16 FILLER_0_61_520 ();
 FILLCELL_X1 FILLER_0_61_536 ();
 FILLCELL_X32 FILLER_0_61_1008 ();
 FILLCELL_X4 FILLER_0_61_1040 ();
 FILLCELL_X2 FILLER_0_61_1044 ();
 FILLCELL_X32 FILLER_0_62_1 ();
 FILLCELL_X4 FILLER_0_62_33 ();
 FILLCELL_X32 FILLER_0_62_456 ();
 FILLCELL_X16 FILLER_0_62_488 ();
 FILLCELL_X4 FILLER_0_62_504 ();
 FILLCELL_X16 FILLER_0_62_521 ();
 FILLCELL_X32 FILLER_0_62_1008 ();
 FILLCELL_X4 FILLER_0_62_1040 ();
 FILLCELL_X2 FILLER_0_62_1044 ();
 FILLCELL_X32 FILLER_0_63_1 ();
 FILLCELL_X4 FILLER_0_63_33 ();
 FILLCELL_X32 FILLER_0_63_456 ();
 FILLCELL_X32 FILLER_0_63_488 ();
 FILLCELL_X16 FILLER_0_63_520 ();
 FILLCELL_X1 FILLER_0_63_536 ();
 FILLCELL_X32 FILLER_0_63_1008 ();
 FILLCELL_X4 FILLER_0_63_1040 ();
 FILLCELL_X2 FILLER_0_63_1044 ();
 FILLCELL_X32 FILLER_0_64_1 ();
 FILLCELL_X4 FILLER_0_64_33 ();
 FILLCELL_X32 FILLER_0_64_456 ();
 FILLCELL_X32 FILLER_0_64_488 ();
 FILLCELL_X16 FILLER_0_64_520 ();
 FILLCELL_X1 FILLER_0_64_536 ();
 FILLCELL_X32 FILLER_0_64_1008 ();
 FILLCELL_X4 FILLER_0_64_1040 ();
 FILLCELL_X2 FILLER_0_64_1044 ();
 FILLCELL_X32 FILLER_0_65_1 ();
 FILLCELL_X32 FILLER_0_65_33 ();
 FILLCELL_X16 FILLER_0_65_65 ();
 FILLCELL_X8 FILLER_0_65_81 ();
 FILLCELL_X32 FILLER_0_65_90 ();
 FILLCELL_X32 FILLER_0_65_122 ();
 FILLCELL_X16 FILLER_0_65_154 ();
 FILLCELL_X8 FILLER_0_65_170 ();
 FILLCELL_X32 FILLER_0_65_179 ();
 FILLCELL_X32 FILLER_0_65_211 ();
 FILLCELL_X16 FILLER_0_65_243 ();
 FILLCELL_X8 FILLER_0_65_259 ();
 FILLCELL_X32 FILLER_0_65_268 ();
 FILLCELL_X32 FILLER_0_65_300 ();
 FILLCELL_X16 FILLER_0_65_332 ();
 FILLCELL_X8 FILLER_0_65_348 ();
 FILLCELL_X32 FILLER_0_65_357 ();
 FILLCELL_X32 FILLER_0_65_389 ();
 FILLCELL_X16 FILLER_0_65_421 ();
 FILLCELL_X8 FILLER_0_65_437 ();
 FILLCELL_X32 FILLER_0_65_446 ();
 FILLCELL_X32 FILLER_0_65_478 ();
 FILLCELL_X16 FILLER_0_65_510 ();
 FILLCELL_X8 FILLER_0_65_526 ();
 FILLCELL_X2 FILLER_0_65_535 ();
 FILLCELL_X32 FILLER_0_65_1008 ();
 FILLCELL_X4 FILLER_0_65_1040 ();
 FILLCELL_X2 FILLER_0_65_1044 ();
 FILLCELL_X32 FILLER_0_66_1 ();
 FILLCELL_X32 FILLER_0_66_33 ();
 FILLCELL_X16 FILLER_0_66_65 ();
 FILLCELL_X8 FILLER_0_66_81 ();
 FILLCELL_X32 FILLER_0_66_90 ();
 FILLCELL_X32 FILLER_0_66_122 ();
 FILLCELL_X32 FILLER_0_66_154 ();
 FILLCELL_X32 FILLER_0_66_186 ();
 FILLCELL_X32 FILLER_0_66_218 ();
 FILLCELL_X16 FILLER_0_66_250 ();
 FILLCELL_X1 FILLER_0_66_266 ();
 FILLCELL_X32 FILLER_0_66_268 ();
 FILLCELL_X32 FILLER_0_66_300 ();
 FILLCELL_X32 FILLER_0_66_332 ();
 FILLCELL_X32 FILLER_0_66_364 ();
 FILLCELL_X32 FILLER_0_66_396 ();
 FILLCELL_X16 FILLER_0_66_428 ();
 FILLCELL_X1 FILLER_0_66_444 ();
 FILLCELL_X32 FILLER_0_66_446 ();
 FILLCELL_X32 FILLER_0_66_478 ();
 FILLCELL_X16 FILLER_0_66_510 ();
 FILLCELL_X8 FILLER_0_66_526 ();
 FILLCELL_X2 FILLER_0_66_534 ();
 FILLCELL_X1 FILLER_0_66_536 ();
 FILLCELL_X32 FILLER_0_66_1008 ();
 FILLCELL_X4 FILLER_0_66_1040 ();
 FILLCELL_X2 FILLER_0_66_1044 ();
 FILLCELL_X32 FILLER_0_67_1 ();
 FILLCELL_X32 FILLER_0_67_33 ();
 FILLCELL_X32 FILLER_0_67_65 ();
 FILLCELL_X32 FILLER_0_67_97 ();
 FILLCELL_X32 FILLER_0_67_129 ();
 FILLCELL_X16 FILLER_0_67_161 ();
 FILLCELL_X1 FILLER_0_67_177 ();
 FILLCELL_X32 FILLER_0_67_179 ();
 FILLCELL_X32 FILLER_0_67_211 ();
 FILLCELL_X32 FILLER_0_67_243 ();
 FILLCELL_X32 FILLER_0_67_275 ();
 FILLCELL_X32 FILLER_0_67_307 ();
 FILLCELL_X16 FILLER_0_67_339 ();
 FILLCELL_X1 FILLER_0_67_355 ();
 FILLCELL_X32 FILLER_0_67_357 ();
 FILLCELL_X32 FILLER_0_67_389 ();
 FILLCELL_X32 FILLER_0_67_421 ();
 FILLCELL_X32 FILLER_0_67_453 ();
 FILLCELL_X32 FILLER_0_67_485 ();
 FILLCELL_X16 FILLER_0_67_517 ();
 FILLCELL_X1 FILLER_0_67_533 ();
 FILLCELL_X2 FILLER_0_67_535 ();
 FILLCELL_X32 FILLER_0_67_1008 ();
 FILLCELL_X4 FILLER_0_67_1040 ();
 FILLCELL_X2 FILLER_0_67_1044 ();
 FILLCELL_X32 FILLER_0_68_1 ();
 FILLCELL_X32 FILLER_0_68_33 ();
 FILLCELL_X16 FILLER_0_68_65 ();
 FILLCELL_X8 FILLER_0_68_81 ();
 FILLCELL_X32 FILLER_0_68_90 ();
 FILLCELL_X32 FILLER_0_68_122 ();
 FILLCELL_X32 FILLER_0_68_154 ();
 FILLCELL_X32 FILLER_0_68_186 ();
 FILLCELL_X32 FILLER_0_68_218 ();
 FILLCELL_X16 FILLER_0_68_250 ();
 FILLCELL_X1 FILLER_0_68_266 ();
 FILLCELL_X32 FILLER_0_68_268 ();
 FILLCELL_X32 FILLER_0_68_300 ();
 FILLCELL_X32 FILLER_0_68_332 ();
 FILLCELL_X32 FILLER_0_68_364 ();
 FILLCELL_X32 FILLER_0_68_396 ();
 FILLCELL_X16 FILLER_0_68_428 ();
 FILLCELL_X1 FILLER_0_68_444 ();
 FILLCELL_X32 FILLER_0_68_446 ();
 FILLCELL_X32 FILLER_0_68_478 ();
 FILLCELL_X16 FILLER_0_68_510 ();
 FILLCELL_X8 FILLER_0_68_526 ();
 FILLCELL_X2 FILLER_0_68_534 ();
 FILLCELL_X1 FILLER_0_68_536 ();
 FILLCELL_X32 FILLER_0_68_1008 ();
 FILLCELL_X4 FILLER_0_68_1040 ();
 FILLCELL_X2 FILLER_0_68_1044 ();
 FILLCELL_X32 FILLER_0_69_1 ();
 FILLCELL_X32 FILLER_0_69_33 ();
 FILLCELL_X16 FILLER_0_69_65 ();
 FILLCELL_X8 FILLER_0_69_81 ();
 FILLCELL_X32 FILLER_0_69_90 ();
 FILLCELL_X32 FILLER_0_69_122 ();
 FILLCELL_X16 FILLER_0_69_154 ();
 FILLCELL_X8 FILLER_0_69_170 ();
 FILLCELL_X32 FILLER_0_69_179 ();
 FILLCELL_X32 FILLER_0_69_211 ();
 FILLCELL_X16 FILLER_0_69_243 ();
 FILLCELL_X8 FILLER_0_69_259 ();
 FILLCELL_X32 FILLER_0_69_268 ();
 FILLCELL_X32 FILLER_0_69_300 ();
 FILLCELL_X16 FILLER_0_69_332 ();
 FILLCELL_X8 FILLER_0_69_348 ();
 FILLCELL_X32 FILLER_0_69_357 ();
 FILLCELL_X32 FILLER_0_69_389 ();
 FILLCELL_X16 FILLER_0_69_421 ();
 FILLCELL_X8 FILLER_0_69_437 ();
 FILLCELL_X32 FILLER_0_69_446 ();
 FILLCELL_X32 FILLER_0_69_478 ();
 FILLCELL_X16 FILLER_0_69_510 ();
 FILLCELL_X8 FILLER_0_69_526 ();
 FILLCELL_X32 FILLER_0_69_535 ();
 FILLCELL_X32 FILLER_0_69_567 ();
 FILLCELL_X16 FILLER_0_69_599 ();
 FILLCELL_X8 FILLER_0_69_615 ();
 FILLCELL_X32 FILLER_0_69_624 ();
 FILLCELL_X32 FILLER_0_69_656 ();
 FILLCELL_X16 FILLER_0_69_688 ();
 FILLCELL_X8 FILLER_0_69_704 ();
 FILLCELL_X32 FILLER_0_69_713 ();
 FILLCELL_X16 FILLER_0_69_745 ();
 FILLCELL_X8 FILLER_0_69_761 ();
 FILLCELL_X2 FILLER_0_69_769 ();
 FILLCELL_X1 FILLER_0_69_771 ();
 FILLCELL_X8 FILLER_0_69_785 ();
 FILLCELL_X4 FILLER_0_69_793 ();
 FILLCELL_X1 FILLER_0_69_797 ();
 FILLCELL_X32 FILLER_0_69_802 ();
 FILLCELL_X32 FILLER_0_69_834 ();
 FILLCELL_X16 FILLER_0_69_866 ();
 FILLCELL_X8 FILLER_0_69_882 ();
 FILLCELL_X32 FILLER_0_69_891 ();
 FILLCELL_X32 FILLER_0_69_923 ();
 FILLCELL_X16 FILLER_0_69_955 ();
 FILLCELL_X8 FILLER_0_69_971 ();
 FILLCELL_X32 FILLER_0_69_980 ();
 FILLCELL_X32 FILLER_0_69_1012 ();
 FILLCELL_X2 FILLER_0_69_1044 ();
 FILLCELL_X32 FILLER_0_70_1 ();
 FILLCELL_X32 FILLER_0_70_33 ();
 FILLCELL_X16 FILLER_0_70_65 ();
 FILLCELL_X8 FILLER_0_70_81 ();
 FILLCELL_X32 FILLER_0_70_90 ();
 FILLCELL_X32 FILLER_0_70_122 ();
 FILLCELL_X32 FILLER_0_70_154 ();
 FILLCELL_X32 FILLER_0_70_186 ();
 FILLCELL_X32 FILLER_0_70_218 ();
 FILLCELL_X16 FILLER_0_70_250 ();
 FILLCELL_X1 FILLER_0_70_266 ();
 FILLCELL_X32 FILLER_0_70_268 ();
 FILLCELL_X32 FILLER_0_70_300 ();
 FILLCELL_X32 FILLER_0_70_332 ();
 FILLCELL_X32 FILLER_0_70_364 ();
 FILLCELL_X32 FILLER_0_70_396 ();
 FILLCELL_X16 FILLER_0_70_428 ();
 FILLCELL_X1 FILLER_0_70_444 ();
 FILLCELL_X32 FILLER_0_70_446 ();
 FILLCELL_X32 FILLER_0_70_478 ();
 FILLCELL_X32 FILLER_0_70_510 ();
 FILLCELL_X32 FILLER_0_70_542 ();
 FILLCELL_X32 FILLER_0_70_574 ();
 FILLCELL_X16 FILLER_0_70_606 ();
 FILLCELL_X1 FILLER_0_70_622 ();
 FILLCELL_X32 FILLER_0_70_624 ();
 FILLCELL_X32 FILLER_0_70_656 ();
 FILLCELL_X32 FILLER_0_70_688 ();
 FILLCELL_X32 FILLER_0_70_720 ();
 FILLCELL_X32 FILLER_0_70_752 ();
 FILLCELL_X16 FILLER_0_70_784 ();
 FILLCELL_X1 FILLER_0_70_800 ();
 FILLCELL_X32 FILLER_0_70_802 ();
 FILLCELL_X32 FILLER_0_70_834 ();
 FILLCELL_X32 FILLER_0_70_866 ();
 FILLCELL_X32 FILLER_0_70_898 ();
 FILLCELL_X32 FILLER_0_70_930 ();
 FILLCELL_X16 FILLER_0_70_962 ();
 FILLCELL_X1 FILLER_0_70_978 ();
 FILLCELL_X32 FILLER_0_70_980 ();
 FILLCELL_X32 FILLER_0_70_1012 ();
 FILLCELL_X2 FILLER_0_70_1044 ();
 FILLCELL_X32 FILLER_0_71_1 ();
 FILLCELL_X32 FILLER_0_71_33 ();
 FILLCELL_X32 FILLER_0_71_65 ();
 FILLCELL_X32 FILLER_0_71_97 ();
 FILLCELL_X32 FILLER_0_71_129 ();
 FILLCELL_X16 FILLER_0_71_161 ();
 FILLCELL_X1 FILLER_0_71_177 ();
 FILLCELL_X32 FILLER_0_71_179 ();
 FILLCELL_X32 FILLER_0_71_211 ();
 FILLCELL_X32 FILLER_0_71_243 ();
 FILLCELL_X32 FILLER_0_71_275 ();
 FILLCELL_X32 FILLER_0_71_307 ();
 FILLCELL_X16 FILLER_0_71_339 ();
 FILLCELL_X1 FILLER_0_71_355 ();
 FILLCELL_X32 FILLER_0_71_357 ();
 FILLCELL_X32 FILLER_0_71_389 ();
 FILLCELL_X32 FILLER_0_71_421 ();
 FILLCELL_X32 FILLER_0_71_453 ();
 FILLCELL_X32 FILLER_0_71_485 ();
 FILLCELL_X16 FILLER_0_71_517 ();
 FILLCELL_X1 FILLER_0_71_533 ();
 FILLCELL_X32 FILLER_0_71_535 ();
 FILLCELL_X32 FILLER_0_71_567 ();
 FILLCELL_X32 FILLER_0_71_599 ();
 FILLCELL_X32 FILLER_0_71_631 ();
 FILLCELL_X32 FILLER_0_71_663 ();
 FILLCELL_X16 FILLER_0_71_695 ();
 FILLCELL_X1 FILLER_0_71_711 ();
 FILLCELL_X32 FILLER_0_71_713 ();
 FILLCELL_X32 FILLER_0_71_745 ();
 FILLCELL_X32 FILLER_0_71_777 ();
 FILLCELL_X32 FILLER_0_71_809 ();
 FILLCELL_X32 FILLER_0_71_841 ();
 FILLCELL_X16 FILLER_0_71_873 ();
 FILLCELL_X1 FILLER_0_71_889 ();
 FILLCELL_X32 FILLER_0_71_891 ();
 FILLCELL_X32 FILLER_0_71_923 ();
 FILLCELL_X32 FILLER_0_71_955 ();
 FILLCELL_X32 FILLER_0_71_987 ();
 FILLCELL_X16 FILLER_0_71_1019 ();
 FILLCELL_X8 FILLER_0_71_1035 ();
 FILLCELL_X2 FILLER_0_71_1043 ();
 FILLCELL_X1 FILLER_0_71_1045 ();
 FILLCELL_X32 FILLER_0_72_1 ();
 FILLCELL_X32 FILLER_0_72_33 ();
 FILLCELL_X16 FILLER_0_72_65 ();
 FILLCELL_X8 FILLER_0_72_81 ();
 FILLCELL_X32 FILLER_0_72_90 ();
 FILLCELL_X32 FILLER_0_72_122 ();
 FILLCELL_X16 FILLER_0_72_154 ();
 FILLCELL_X8 FILLER_0_72_170 ();
 FILLCELL_X32 FILLER_0_72_179 ();
 FILLCELL_X32 FILLER_0_72_211 ();
 FILLCELL_X4 FILLER_0_72_243 ();
 FILLCELL_X2 FILLER_0_72_247 ();
 FILLCELL_X1 FILLER_0_72_249 ();
 FILLCELL_X8 FILLER_0_72_252 ();
 FILLCELL_X4 FILLER_0_72_260 ();
 FILLCELL_X2 FILLER_0_72_264 ();
 FILLCELL_X1 FILLER_0_72_266 ();
 FILLCELL_X32 FILLER_0_72_268 ();
 FILLCELL_X32 FILLER_0_72_300 ();
 FILLCELL_X16 FILLER_0_72_332 ();
 FILLCELL_X8 FILLER_0_72_348 ();
 FILLCELL_X32 FILLER_0_72_357 ();
 FILLCELL_X32 FILLER_0_72_389 ();
 FILLCELL_X16 FILLER_0_72_421 ();
 FILLCELL_X8 FILLER_0_72_437 ();
 FILLCELL_X32 FILLER_0_72_446 ();
 FILLCELL_X32 FILLER_0_72_478 ();
 FILLCELL_X16 FILLER_0_72_510 ();
 FILLCELL_X8 FILLER_0_72_526 ();
 FILLCELL_X32 FILLER_0_72_535 ();
 FILLCELL_X32 FILLER_0_72_567 ();
 FILLCELL_X16 FILLER_0_72_599 ();
 FILLCELL_X8 FILLER_0_72_615 ();
 FILLCELL_X32 FILLER_0_72_624 ();
 FILLCELL_X32 FILLER_0_72_656 ();
 FILLCELL_X16 FILLER_0_72_688 ();
 FILLCELL_X8 FILLER_0_72_704 ();
 FILLCELL_X32 FILLER_0_72_713 ();
 FILLCELL_X32 FILLER_0_72_745 ();
 FILLCELL_X16 FILLER_0_72_777 ();
 FILLCELL_X8 FILLER_0_72_793 ();
 FILLCELL_X32 FILLER_0_72_802 ();
 FILLCELL_X32 FILLER_0_72_834 ();
 FILLCELL_X16 FILLER_0_72_866 ();
 FILLCELL_X8 FILLER_0_72_882 ();
 FILLCELL_X32 FILLER_0_72_891 ();
 FILLCELL_X32 FILLER_0_72_923 ();
 FILLCELL_X16 FILLER_0_72_955 ();
 FILLCELL_X8 FILLER_0_72_971 ();
 FILLCELL_X32 FILLER_0_72_980 ();
 FILLCELL_X32 FILLER_0_72_1012 ();
 FILLCELL_X2 FILLER_0_72_1044 ();
endmodule
