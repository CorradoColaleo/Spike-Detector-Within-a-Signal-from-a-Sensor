module iir (clk,
    rst,
    x,
    z);
 input clk;
 input rst;
 input [10:0] x;
 output [10:0] z;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire \iir1.t1[0] ;
 wire \iir1.t1[1] ;
 wire \iir1.t1[2] ;
 wire \iir1.t1[3] ;
 wire \iir1.t1[4] ;
 wire \iir1.x1[10] ;
 wire \iir1.x1[5] ;
 wire \iir1.x1[6] ;
 wire \iir1.x1[7] ;
 wire \iir1.x1[8] ;
 wire \iir1.x1[9] ;
 wire \iir1.x2[0] ;
 wire \iir1.x2[10] ;
 wire \iir1.x2[1] ;
 wire \iir1.x2[2] ;
 wire \iir1.x2[3] ;
 wire \iir1.x2[4] ;
 wire \iir1.x2[5] ;
 wire \iir1.x2[6] ;
 wire \iir1.x2[7] ;
 wire \iir1.x2[8] ;
 wire \iir1.x2[9] ;
 wire \iir1.x[0] ;
 wire \iir1.x[10] ;
 wire \iir1.x[1] ;
 wire \iir1.x[2] ;
 wire \iir1.x[3] ;
 wire \iir1.x[4] ;
 wire \iir1.x[5] ;
 wire \iir1.x[6] ;
 wire \iir1.x[7] ;
 wire \iir1.x[8] ;
 wire \iir1.x[9] ;
 wire \iir1.y2[0] ;
 wire \iir1.y2[10] ;
 wire \iir1.y2[1] ;
 wire \iir1.y2[2] ;
 wire \iir1.y2[3] ;
 wire \iir1.y2[4] ;
 wire \iir1.y2[5] ;
 wire \iir1.y2[6] ;
 wire \iir1.y2[7] ;
 wire \iir1.y2[8] ;
 wire \iir1.y2[9] ;
 wire \iir1.y[0] ;
 wire \iir1.y[10] ;
 wire \iir1.y[1] ;
 wire \iir1.y[2] ;
 wire \iir1.y[3] ;
 wire \iir1.y[4] ;
 wire \iir1.y[5] ;
 wire \iir1.y[6] ;
 wire \iir1.y[7] ;
 wire \iir1.y[8] ;
 wire \iir1.y[9] ;
 wire \iir2.x2[0] ;
 wire \iir2.x2[10] ;
 wire \iir2.x2[1] ;
 wire \iir2.x2[2] ;
 wire \iir2.x2[3] ;
 wire \iir2.x2[4] ;
 wire \iir2.x2[5] ;
 wire \iir2.x2[6] ;
 wire \iir2.x2[7] ;
 wire \iir2.x2[8] ;
 wire \iir2.x2[9] ;
 wire \iir2.y2[0] ;
 wire \iir2.y2[10] ;
 wire \iir2.y2[1] ;
 wire \iir2.y2[2] ;
 wire \iir2.y2[3] ;
 wire \iir2.y2[4] ;
 wire \iir2.y2[5] ;
 wire \iir2.y2[6] ;
 wire \iir2.y2[7] ;
 wire \iir2.y2[8] ;
 wire \iir2.y2[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;

 INV_X1 _3008_ (.A(rst),
    .ZN(_1297_));
 XNOR2_X1 _3009_ (.A(\iir2.y2[10] ),
    .B(\iir2.y2[8] ),
    .ZN(_1308_));
 INV_X1 _3010_ (.A(_1308_),
    .ZN(_1319_));
 XNOR2_X1 _3011_ (.A(z[1]),
    .B(z[0]),
    .ZN(_1330_));
 INV_X1 _3012_ (.A(\iir2.x2[4] ),
    .ZN(_1341_));
 NOR3_X1 _3013_ (.A1(\iir1.y[2] ),
    .A2(\iir1.y[1] ),
    .A3(\iir1.y[0] ),
    .ZN(_1352_));
 XOR2_X1 _3014_ (.A(\iir1.y[3] ),
    .B(_1352_),
    .Z(_1363_));
 XNOR2_X1 _3015_ (.A(\iir1.y2[2] ),
    .B(_1363_),
    .ZN(_1374_));
 XOR2_X1 _3016_ (.A(\iir1.y[1] ),
    .B(\iir1.y[0] ),
    .Z(_1385_));
 NAND2_X1 _3017_ (.A1(\iir1.y2[0] ),
    .A2(_1385_),
    .ZN(_1396_));
 INV_X1 _3018_ (.A(net84),
    .ZN(_1407_));
 NAND2_X1 _3019_ (.A1(\iir1.y[2] ),
    .A2(\iir1.y[1] ),
    .ZN(_1418_));
 XOR2_X1 _3020_ (.A(\iir1.y[2] ),
    .B(\iir1.y[0] ),
    .Z(_1429_));
 OR2_X1 _3021_ (.A1(\iir1.y[1] ),
    .A2(_1429_),
    .ZN(_1440_));
 NAND2_X1 _3022_ (.A1(_1418_),
    .A2(_1440_),
    .ZN(_1451_));
 XNOR2_X1 _3023_ (.A(_1407_),
    .B(_1451_),
    .ZN(_1462_));
 NOR2_X1 _3024_ (.A1(_1396_),
    .A2(_1462_),
    .ZN(_1473_));
 NAND2_X1 _3025_ (.A1(_1374_),
    .A2(_1473_),
    .ZN(_1484_));
 NAND4_X1 _3026_ (.A1(\iir1.y2[1] ),
    .A2(_1418_),
    .A3(_1374_),
    .A4(_1440_),
    .ZN(_1495_));
 INV_X1 _3027_ (.A(net76),
    .ZN(_1506_));
 OR2_X1 _3028_ (.A1(_1506_),
    .A2(_1363_),
    .ZN(_1517_));
 AND3_X1 _3029_ (.A1(\iir1.y[3] ),
    .A2(\iir1.y[2] ),
    .A3(\iir1.y[1] ),
    .ZN(_1528_));
 NAND2_X1 _3030_ (.A1(\iir1.y[0] ),
    .A2(_1528_),
    .ZN(_1539_));
 XOR2_X1 _3031_ (.A(\iir1.y[4] ),
    .B(\iir1.y[3] ),
    .Z(_1550_));
 XNOR2_X1 _3032_ (.A(\iir1.y[2] ),
    .B(_1550_),
    .ZN(_1561_));
 NAND2_X1 _3033_ (.A1(\iir1.y[3] ),
    .A2(\iir1.y[2] ),
    .ZN(_1572_));
 OAI21_X1 _3034_ (.A(\iir1.y[1] ),
    .B1(\iir1.y[2] ),
    .B2(\iir1.y[3] ),
    .ZN(_1583_));
 NAND2_X1 _3035_ (.A1(_1572_),
    .A2(_1583_),
    .ZN(_1594_));
 XNOR2_X1 _3036_ (.A(_1561_),
    .B(_1594_),
    .ZN(_1605_));
 XNOR2_X1 _3037_ (.A(\iir1.y[1] ),
    .B(_1605_),
    .ZN(_1616_));
 OR2_X1 _3038_ (.A1(\iir1.y[3] ),
    .A2(\iir1.y[2] ),
    .ZN(_1627_));
 OAI22_X1 _3039_ (.A1(\iir1.y[0] ),
    .A2(_1528_),
    .B1(_1627_),
    .B2(\iir1.y[1] ),
    .ZN(_1638_));
 XOR2_X1 _3040_ (.A(_1616_),
    .B(_1638_),
    .Z(_1649_));
 XNOR2_X1 _3041_ (.A(_1539_),
    .B(_1649_),
    .ZN(_1660_));
 XNOR2_X1 _3042_ (.A(_0012_),
    .B(_1660_),
    .ZN(_1671_));
 XOR2_X1 _3043_ (.A(_1517_),
    .B(_1671_),
    .Z(_1682_));
 XNOR2_X1 _3044_ (.A(_0015_),
    .B(_1682_),
    .ZN(_1693_));
 XNOR2_X1 _3045_ (.A(_1495_),
    .B(_1693_),
    .ZN(_1704_));
 XNOR2_X1 _3046_ (.A(_1484_),
    .B(_1704_),
    .ZN(_1715_));
 XNOR2_X1 _3047_ (.A(_1341_),
    .B(_1715_),
    .ZN(_1726_));
 XNOR2_X1 _3048_ (.A(\iir2.x2[3] ),
    .B(_1726_),
    .ZN(_1737_));
 OAI22_X1 _3049_ (.A1(_1407_),
    .A2(_1451_),
    .B1(_1396_),
    .B2(_1462_),
    .ZN(_1748_));
 XNOR2_X1 _3050_ (.A(_1374_),
    .B(_1748_),
    .ZN(_1759_));
 NOR2_X1 _3051_ (.A1(_0021_),
    .A2(_1759_),
    .ZN(_1770_));
 XNOR2_X1 _3052_ (.A(\iir2.x2[3] ),
    .B(_1759_),
    .ZN(_1781_));
 AND2_X1 _3053_ (.A1(\iir2.x2[2] ),
    .A2(_1781_),
    .ZN(_1792_));
 OAI21_X1 _3054_ (.A(_1737_),
    .B1(_1770_),
    .B2(_1792_),
    .ZN(_1803_));
 OR3_X1 _3055_ (.A1(_1792_),
    .A2(_1770_),
    .A3(_1737_),
    .ZN(_1814_));
 AND2_X1 _3056_ (.A1(_1803_),
    .A2(_1814_),
    .ZN(_1825_));
 XOR2_X1 _3057_ (.A(\iir2.x2[1] ),
    .B(\iir2.x2[2] ),
    .Z(_1836_));
 NAND2_X1 _3058_ (.A1(_1825_),
    .A2(_1836_),
    .ZN(_1847_));
 NAND2_X1 _3059_ (.A1(_1803_),
    .A2(_1847_),
    .ZN(_1858_));
 INV_X1 _3060_ (.A(\iir2.x2[3] ),
    .ZN(_1869_));
 OAI22_X1 _3061_ (.A1(_0019_),
    .A2(_1715_),
    .B1(_1726_),
    .B2(_1869_),
    .ZN(_1880_));
 NOR2_X1 _3062_ (.A1(\iir1.y2[3] ),
    .A2(_1660_),
    .ZN(_1891_));
 NAND3_X1 _3063_ (.A1(\iir1.y[0] ),
    .A2(_1528_),
    .A3(_1616_),
    .ZN(_1902_));
 NOR2_X1 _3064_ (.A1(_1616_),
    .A2(_1638_),
    .ZN(_1913_));
 AOI21_X1 _3065_ (.A(_1561_),
    .B1(_1583_),
    .B2(_1572_),
    .ZN(_1924_));
 AOI21_X1 _3066_ (.A(_1924_),
    .B1(_1605_),
    .B2(\iir1.y[1] ),
    .ZN(_1935_));
 AND2_X1 _3067_ (.A1(\iir1.y[4] ),
    .A2(\iir1.y[3] ),
    .ZN(_1946_));
 AOI21_X1 _3068_ (.A(_1946_),
    .B1(_1550_),
    .B2(\iir1.y[2] ),
    .ZN(_1957_));
 XOR2_X1 _3069_ (.A(\iir1.y[5] ),
    .B(\iir1.y[3] ),
    .Z(_1968_));
 XNOR2_X1 _3070_ (.A(\iir1.y[4] ),
    .B(_1968_),
    .ZN(_1979_));
 XOR2_X1 _3071_ (.A(_1957_),
    .B(_1979_),
    .Z(_1990_));
 XNOR2_X1 _3072_ (.A(_1429_),
    .B(_1990_),
    .ZN(_2001_));
 XOR2_X1 _3073_ (.A(_1935_),
    .B(_2001_),
    .Z(_2012_));
 XOR2_X1 _3074_ (.A(_1913_),
    .B(_2012_),
    .Z(_2023_));
 XNOR2_X1 _3075_ (.A(_1902_),
    .B(_2023_),
    .ZN(_2034_));
 XNOR2_X1 _3076_ (.A(_0011_),
    .B(_2034_),
    .ZN(_2045_));
 XNOR2_X1 _3077_ (.A(_1891_),
    .B(_2045_),
    .ZN(_2056_));
 XNOR2_X1 _3078_ (.A(_0014_),
    .B(_2056_),
    .ZN(_2067_));
 NAND2_X1 _3079_ (.A1(_0015_),
    .A2(_1682_),
    .ZN(_2078_));
 OR2_X1 _3080_ (.A1(_1517_),
    .A2(_1671_),
    .ZN(_2089_));
 AOI21_X1 _3081_ (.A(_2067_),
    .B1(_2078_),
    .B2(_2089_),
    .ZN(_2100_));
 AND3_X1 _3082_ (.A1(_2089_),
    .A2(_2078_),
    .A3(_2067_),
    .ZN(_2111_));
 NOR2_X1 _3083_ (.A1(_2100_),
    .A2(_2111_),
    .ZN(_2122_));
 OR2_X1 _3084_ (.A1(_1495_),
    .A2(_1693_),
    .ZN(_2133_));
 OAI21_X1 _3085_ (.A(_2133_),
    .B1(_1704_),
    .B2(_1484_),
    .ZN(_2144_));
 XNOR2_X1 _3086_ (.A(_2122_),
    .B(_2144_),
    .ZN(_2155_));
 XOR2_X1 _3087_ (.A(\iir2.x2[5] ),
    .B(_2155_),
    .Z(_2166_));
 XNOR2_X1 _3088_ (.A(\iir2.x2[4] ),
    .B(_2166_),
    .ZN(_2177_));
 XNOR2_X1 _3089_ (.A(_1880_),
    .B(_2177_),
    .ZN(_2188_));
 XNOR2_X1 _3090_ (.A(\iir2.x2[2] ),
    .B(\iir2.x2[3] ),
    .ZN(_2199_));
 XOR2_X1 _3091_ (.A(_2188_),
    .B(_2199_),
    .Z(_2210_));
 AND2_X1 _3092_ (.A1(_1858_),
    .A2(_2210_),
    .ZN(_2221_));
 XOR2_X1 _3093_ (.A(_1858_),
    .B(_2210_),
    .Z(_2229_));
 NAND2_X1 _3094_ (.A1(\iir2.x2[1] ),
    .A2(\iir2.x2[2] ),
    .ZN(_2235_));
 XOR2_X1 _3095_ (.A(_0024_),
    .B(_2235_),
    .Z(_2245_));
 AOI21_X1 _3096_ (.A(_2221_),
    .B1(_2229_),
    .B2(_2245_),
    .ZN(_2256_));
 NAND2_X1 _3097_ (.A1(_1880_),
    .A2(_2177_),
    .ZN(_2262_));
 OAI21_X1 _3098_ (.A(_2262_),
    .B1(_2188_),
    .B2(_2199_),
    .ZN(_2263_));
 OAI22_X1 _3099_ (.A1(_0017_),
    .A2(_2155_),
    .B1(_2166_),
    .B2(_1341_),
    .ZN(_2264_));
 INV_X1 _3100_ (.A(\iir2.x2[6] ),
    .ZN(_2265_));
 OAI21_X1 _3101_ (.A(_2045_),
    .B1(_1660_),
    .B2(\iir1.y2[3] ),
    .ZN(_2266_));
 NAND2_X1 _3102_ (.A1(_0014_),
    .A2(_2056_),
    .ZN(_2267_));
 NAND2_X1 _3103_ (.A1(_2266_),
    .A2(_2267_),
    .ZN(_2268_));
 NAND2_X1 _3104_ (.A1(\iir1.y2[4] ),
    .A2(_2034_),
    .ZN(_2269_));
 NAND4_X1 _3105_ (.A1(\iir1.y[0] ),
    .A2(_1528_),
    .A3(_1616_),
    .A4(_2012_),
    .ZN(_2270_));
 AND2_X1 _3106_ (.A1(\iir1.y[2] ),
    .A2(\iir1.y[0] ),
    .ZN(_2271_));
 NOR2_X1 _3107_ (.A1(_1957_),
    .A2(_1979_),
    .ZN(_2272_));
 AOI21_X1 _3108_ (.A(_2272_),
    .B1(_1990_),
    .B2(_1429_),
    .ZN(_2273_));
 XOR2_X1 _3109_ (.A(\iir1.y[3] ),
    .B(\iir1.y[1] ),
    .Z(_2274_));
 NOR2_X1 _3110_ (.A1(\iir1.y[4] ),
    .A2(\iir1.y[3] ),
    .ZN(_2275_));
 NAND2_X1 _3111_ (.A1(\iir1.y[4] ),
    .A2(\iir1.y[3] ),
    .ZN(_2276_));
 INV_X1 _3112_ (.A(net86),
    .ZN(_2277_));
 AOI21_X1 _3113_ (.A(_2275_),
    .B1(_2276_),
    .B2(_2277_),
    .ZN(_2278_));
 XOR2_X1 _3114_ (.A(\iir1.y[6] ),
    .B(\iir1.y[5] ),
    .Z(_2279_));
 XNOR2_X1 _3115_ (.A(\iir1.y[4] ),
    .B(_2279_),
    .ZN(_2280_));
 XNOR2_X1 _3116_ (.A(_2278_),
    .B(_2280_),
    .ZN(_2281_));
 XNOR2_X1 _3117_ (.A(_2274_),
    .B(_2281_),
    .ZN(_2282_));
 XOR2_X1 _3118_ (.A(_2273_),
    .B(_2282_),
    .Z(_2283_));
 XOR2_X1 _3119_ (.A(_2271_),
    .B(_2283_),
    .Z(_2284_));
 NOR2_X1 _3120_ (.A1(_1935_),
    .A2(_2001_),
    .ZN(_2285_));
 AOI21_X1 _3121_ (.A(_2285_),
    .B1(_2012_),
    .B2(_1913_),
    .ZN(_2286_));
 XOR2_X1 _3122_ (.A(_2284_),
    .B(_2286_),
    .Z(_2287_));
 XOR2_X1 _3123_ (.A(_2270_),
    .B(_2287_),
    .Z(_2288_));
 XNOR2_X1 _3124_ (.A(\iir1.y2[5] ),
    .B(_2288_),
    .ZN(_2289_));
 XOR2_X1 _3125_ (.A(_2269_),
    .B(_2289_),
    .Z(_2290_));
 XNOR2_X1 _3126_ (.A(\iir1.y2[2] ),
    .B(_2290_),
    .ZN(_2291_));
 XOR2_X1 _3127_ (.A(_2268_),
    .B(_2291_),
    .Z(_2292_));
 AOI21_X1 _3128_ (.A(_2100_),
    .B1(_2122_),
    .B2(_2144_),
    .ZN(_2293_));
 XNOR2_X1 _3129_ (.A(_2292_),
    .B(_2293_),
    .ZN(_2294_));
 XNOR2_X1 _3130_ (.A(_2265_),
    .B(_2294_),
    .ZN(_2295_));
 XOR2_X1 _3131_ (.A(\iir2.x2[5] ),
    .B(_2295_),
    .Z(_2296_));
 XNOR2_X1 _3132_ (.A(_2264_),
    .B(_2296_),
    .ZN(_2297_));
 XNOR2_X1 _3133_ (.A(\iir2.x2[3] ),
    .B(\iir2.x2[4] ),
    .ZN(_2298_));
 XOR2_X1 _3134_ (.A(_2297_),
    .B(_2298_),
    .Z(_2299_));
 XNOR2_X1 _3135_ (.A(_2263_),
    .B(_2299_),
    .ZN(_2300_));
 NAND2_X1 _3136_ (.A1(\iir2.x2[2] ),
    .A2(\iir2.x2[3] ),
    .ZN(_2301_));
 XOR2_X1 _3137_ (.A(_0023_),
    .B(_2301_),
    .Z(_2302_));
 XNOR2_X1 _3138_ (.A(_2300_),
    .B(_2302_),
    .ZN(_2303_));
 INV_X1 _3139_ (.A(_2303_),
    .ZN(_2304_));
 NOR2_X1 _3140_ (.A1(_2256_),
    .A2(_2304_),
    .ZN(_2305_));
 XNOR2_X1 _3141_ (.A(_2256_),
    .B(_2303_),
    .ZN(_2306_));
 NOR2_X1 _3142_ (.A1(_0024_),
    .A2(_2235_),
    .ZN(_2307_));
 AOI21_X1 _3143_ (.A(_2305_),
    .B1(_2306_),
    .B2(_2307_),
    .ZN(_2308_));
 OR2_X1 _3144_ (.A1(_0023_),
    .A2(_2301_),
    .ZN(_2309_));
 NAND2_X1 _3145_ (.A1(_2263_),
    .A2(_2299_),
    .ZN(_2310_));
 INV_X1 _3146_ (.A(_2302_),
    .ZN(_2311_));
 OAI21_X1 _3147_ (.A(_2310_),
    .B1(_2300_),
    .B2(_2311_),
    .ZN(_2312_));
 NAND2_X1 _3148_ (.A1(_2264_),
    .A2(_2296_),
    .ZN(_2313_));
 OAI21_X1 _3149_ (.A(_2313_),
    .B1(_2297_),
    .B2(_2298_),
    .ZN(_2314_));
 AND2_X1 _3150_ (.A1(\iir2.x2[5] ),
    .A2(_2295_),
    .ZN(_2315_));
 INV_X1 _3151_ (.A(_0020_),
    .ZN(_2316_));
 AND2_X1 _3152_ (.A1(_2316_),
    .A2(_2294_),
    .ZN(_2317_));
 NOR2_X1 _3153_ (.A1(_2315_),
    .A2(_2317_),
    .ZN(_2318_));
 INV_X1 _3154_ (.A(\iir2.x2[7] ),
    .ZN(_2319_));
 NAND2_X1 _3155_ (.A1(_2268_),
    .A2(_2291_),
    .ZN(_2320_));
 NAND2_X1 _3156_ (.A1(\iir1.y2[5] ),
    .A2(_2288_),
    .ZN(_2321_));
 NAND3_X1 _3157_ (.A1(_1913_),
    .A2(_2012_),
    .A3(_2284_),
    .ZN(_2322_));
 OAI21_X1 _3158_ (.A(_2322_),
    .B1(_2287_),
    .B2(_2270_),
    .ZN(_2323_));
 NAND2_X1 _3159_ (.A1(_2285_),
    .A2(_2284_),
    .ZN(_2324_));
 NOR2_X1 _3160_ (.A1(_2273_),
    .A2(_2282_),
    .ZN(_2325_));
 AOI21_X1 _3161_ (.A(_2325_),
    .B1(_2283_),
    .B2(_2271_),
    .ZN(_2326_));
 NAND2_X1 _3162_ (.A1(\iir1.y[3] ),
    .A2(\iir1.y[1] ),
    .ZN(_2327_));
 INV_X1 _3163_ (.A(_2327_),
    .ZN(_2328_));
 AOI211_X1 _3164_ (.A(_2275_),
    .B(_2280_),
    .C1(_2276_),
    .C2(_2277_),
    .ZN(_2329_));
 AOI21_X1 _3165_ (.A(_2329_),
    .B1(_2281_),
    .B2(_2274_),
    .ZN(_2330_));
 AND2_X1 _3166_ (.A1(\iir1.y[6] ),
    .A2(\iir1.y[5] ),
    .ZN(_2331_));
 AOI21_X1 _3167_ (.A(_2331_),
    .B1(_2279_),
    .B2(\iir1.y[4] ),
    .ZN(_2332_));
 XOR2_X1 _3168_ (.A(\iir1.y[7] ),
    .B(\iir1.y[6] ),
    .Z(_2333_));
 XNOR2_X1 _3169_ (.A(_0007_),
    .B(_2333_),
    .ZN(_2334_));
 XOR2_X1 _3170_ (.A(_2332_),
    .B(_2334_),
    .Z(_2335_));
 XNOR2_X1 _3171_ (.A(\iir1.y[4] ),
    .B(\iir1.y[2] ),
    .ZN(_2336_));
 XNOR2_X1 _3172_ (.A(_2335_),
    .B(_2336_),
    .ZN(_2337_));
 XOR2_X1 _3173_ (.A(_2330_),
    .B(_2337_),
    .Z(_2338_));
 XNOR2_X1 _3174_ (.A(_2328_),
    .B(_2338_),
    .ZN(_2339_));
 XOR2_X1 _3175_ (.A(_2326_),
    .B(_2339_),
    .Z(_2340_));
 XNOR2_X1 _3176_ (.A(_2324_),
    .B(_2340_),
    .ZN(_2341_));
 XNOR2_X1 _3177_ (.A(_2323_),
    .B(_2341_),
    .ZN(_2342_));
 XNOR2_X1 _3178_ (.A(\iir1.y2[6] ),
    .B(_2342_),
    .ZN(_2343_));
 XNOR2_X1 _3179_ (.A(_2321_),
    .B(_2343_),
    .ZN(_2344_));
 XNOR2_X1 _3180_ (.A(\iir1.y2[3] ),
    .B(_2344_),
    .ZN(_2345_));
 NOR2_X1 _3181_ (.A1(_2269_),
    .A2(_2289_),
    .ZN(_2346_));
 AOI21_X1 _3182_ (.A(_2346_),
    .B1(_2290_),
    .B2(_0013_),
    .ZN(_2347_));
 XOR2_X1 _3183_ (.A(_2345_),
    .B(_2347_),
    .Z(_2348_));
 XOR2_X1 _3184_ (.A(_2320_),
    .B(_2348_),
    .Z(_2349_));
 INV_X1 _3185_ (.A(_2292_),
    .ZN(_2350_));
 NOR2_X1 _3186_ (.A1(_2350_),
    .A2(_2293_),
    .ZN(_2351_));
 XNOR2_X1 _3187_ (.A(_2349_),
    .B(_2351_),
    .ZN(_2352_));
 XNOR2_X1 _3188_ (.A(_2319_),
    .B(_2352_),
    .ZN(_2353_));
 XNOR2_X1 _3189_ (.A(\iir2.x2[6] ),
    .B(_2353_),
    .ZN(_2354_));
 XNOR2_X1 _3190_ (.A(_2318_),
    .B(_2354_),
    .ZN(_2355_));
 XOR2_X1 _3191_ (.A(\iir2.x2[4] ),
    .B(\iir2.x2[5] ),
    .Z(_2356_));
 XNOR2_X1 _3192_ (.A(_2355_),
    .B(_2356_),
    .ZN(_2357_));
 XOR2_X1 _3193_ (.A(_2314_),
    .B(_2357_),
    .Z(_2358_));
 NAND2_X1 _3194_ (.A1(\iir2.x2[3] ),
    .A2(\iir2.x2[4] ),
    .ZN(_2359_));
 XOR2_X1 _3195_ (.A(_0022_),
    .B(_2359_),
    .Z(_2360_));
 XNOR2_X1 _3196_ (.A(_2358_),
    .B(_2360_),
    .ZN(_2361_));
 XNOR2_X1 _3197_ (.A(_2312_),
    .B(_2361_),
    .ZN(_2362_));
 XNOR2_X1 _3198_ (.A(_2309_),
    .B(_2362_),
    .ZN(_2363_));
 NOR2_X1 _3199_ (.A1(_2308_),
    .A2(_2363_),
    .ZN(_2364_));
 XOR2_X1 _3200_ (.A(_2308_),
    .B(_2363_),
    .Z(_2365_));
 XNOR2_X1 _3201_ (.A(_2229_),
    .B(_2245_),
    .ZN(_2366_));
 NAND2_X1 _3202_ (.A1(\iir2.x2[0] ),
    .A2(\iir2.x2[1] ),
    .ZN(_2367_));
 XNOR2_X1 _3203_ (.A(_1396_),
    .B(_1462_),
    .ZN(_2368_));
 XOR2_X1 _3204_ (.A(\iir2.x2[2] ),
    .B(_2368_),
    .Z(_2369_));
 INV_X1 _3205_ (.A(\iir2.x2[1] ),
    .ZN(_2370_));
 OAI22_X1 _3206_ (.A1(_0022_),
    .A2(_2368_),
    .B1(_2369_),
    .B2(_2370_),
    .ZN(_2371_));
 XOR2_X1 _3207_ (.A(\iir2.x2[2] ),
    .B(_1781_),
    .Z(_2372_));
 NAND2_X1 _3208_ (.A1(_2371_),
    .A2(_2372_),
    .ZN(_2373_));
 XNOR2_X1 _3209_ (.A(\iir2.x2[0] ),
    .B(\iir2.x2[1] ),
    .ZN(_2374_));
 XNOR2_X1 _3210_ (.A(_2371_),
    .B(_2372_),
    .ZN(_2375_));
 OAI21_X1 _3211_ (.A(_2373_),
    .B1(_2374_),
    .B2(_2375_),
    .ZN(_2376_));
 XOR2_X1 _3212_ (.A(_1825_),
    .B(_1836_),
    .Z(_2377_));
 XNOR2_X1 _3213_ (.A(_2376_),
    .B(_2377_),
    .ZN(_2378_));
 OR2_X1 _3214_ (.A1(_2367_),
    .A2(_2378_),
    .ZN(_2379_));
 NAND2_X1 _3215_ (.A1(_2376_),
    .A2(_2377_),
    .ZN(_2380_));
 AOI21_X1 _3216_ (.A(_2366_),
    .B1(_2379_),
    .B2(_2380_),
    .ZN(_2381_));
 XOR2_X1 _3217_ (.A(_2307_),
    .B(_2306_),
    .Z(_2382_));
 NAND2_X1 _3218_ (.A1(_2381_),
    .A2(_2382_),
    .ZN(_2383_));
 XNOR2_X1 _3219_ (.A(_2374_),
    .B(_2375_),
    .ZN(_2384_));
 INV_X1 _3220_ (.A(net47),
    .ZN(_2385_));
 XNOR2_X1 _3221_ (.A(_2385_),
    .B(_1385_),
    .ZN(_2386_));
 INV_X1 _3222_ (.A(_2386_),
    .ZN(_2387_));
 XNOR2_X1 _3223_ (.A(\iir2.x2[1] ),
    .B(_2386_),
    .ZN(_2388_));
 INV_X1 _3224_ (.A(\iir2.x2[0] ),
    .ZN(_2389_));
 OAI22_X1 _3225_ (.A1(_0023_),
    .A2(_2387_),
    .B1(_2388_),
    .B2(_2389_),
    .ZN(_2390_));
 XNOR2_X1 _3226_ (.A(\iir2.x2[1] ),
    .B(_2369_),
    .ZN(_2391_));
 AND2_X1 _3227_ (.A1(_2390_),
    .A2(_2391_),
    .ZN(_2392_));
 XOR2_X1 _3228_ (.A(_2390_),
    .B(_2391_),
    .Z(_2393_));
 AOI21_X1 _3229_ (.A(_2392_),
    .B1(_2393_),
    .B2(\iir2.x2[0] ),
    .ZN(_2394_));
 NOR2_X1 _3230_ (.A1(_2384_),
    .A2(_2394_),
    .ZN(_2395_));
 XOR2_X1 _3231_ (.A(_2367_),
    .B(_2378_),
    .Z(_2396_));
 NAND2_X1 _3232_ (.A1(_2395_),
    .A2(_2396_),
    .ZN(_2397_));
 AND3_X1 _3233_ (.A1(_2380_),
    .A2(_2379_),
    .A3(_2366_),
    .ZN(_2398_));
 OR2_X1 _3234_ (.A1(_2381_),
    .A2(_2398_),
    .ZN(_2399_));
 NOR2_X1 _3235_ (.A1(_2397_),
    .A2(_2399_),
    .ZN(_2400_));
 NAND3_X1 _3236_ (.A1(\iir1.y[0] ),
    .A2(\iir2.x2[0] ),
    .A3(_2388_),
    .ZN(_2401_));
 NOR2_X1 _3237_ (.A1(_2393_),
    .A2(_2401_),
    .ZN(_2402_));
 XOR2_X1 _3238_ (.A(_2384_),
    .B(_2394_),
    .Z(_2403_));
 NAND2_X1 _3239_ (.A1(_2402_),
    .A2(_2403_),
    .ZN(_2404_));
 XNOR2_X1 _3240_ (.A(_2395_),
    .B(_2396_),
    .ZN(_2405_));
 OR2_X1 _3241_ (.A1(_2404_),
    .A2(_2405_),
    .ZN(_2406_));
 INV_X1 _3242_ (.A(_2406_),
    .ZN(_2407_));
 XOR2_X1 _3243_ (.A(_2397_),
    .B(_2399_),
    .Z(_2408_));
 AOI21_X1 _3244_ (.A(_2400_),
    .B1(_2407_),
    .B2(_2408_),
    .ZN(_2409_));
 XNOR2_X1 _3245_ (.A(_2381_),
    .B(_2382_),
    .ZN(_2410_));
 OAI21_X1 _3246_ (.A(_2383_),
    .B1(_2409_),
    .B2(_2410_),
    .ZN(_2411_));
 AOI21_X1 _3247_ (.A(_2364_),
    .B1(_2365_),
    .B2(_2411_),
    .ZN(_2412_));
 NAND2_X1 _3248_ (.A1(_2312_),
    .A2(_2361_),
    .ZN(_2413_));
 OAI21_X1 _3249_ (.A(_2413_),
    .B1(_2362_),
    .B2(_2309_),
    .ZN(_2414_));
 NOR2_X1 _3250_ (.A1(_0022_),
    .A2(_2359_),
    .ZN(_2415_));
 INV_X1 _3251_ (.A(_2357_),
    .ZN(_2416_));
 NAND2_X1 _3252_ (.A1(_2314_),
    .A2(_2416_),
    .ZN(_2417_));
 INV_X1 _3253_ (.A(_2360_),
    .ZN(_2418_));
 OR2_X1 _3254_ (.A1(_2358_),
    .A2(_2418_),
    .ZN(_2419_));
 NAND2_X1 _3255_ (.A1(_2417_),
    .A2(_2419_),
    .ZN(_2420_));
 OAI21_X1 _3256_ (.A(_2354_),
    .B1(_2317_),
    .B2(_2315_),
    .ZN(_2421_));
 NAND2_X1 _3257_ (.A1(_2355_),
    .A2(_2356_),
    .ZN(_2422_));
 NAND2_X1 _3258_ (.A1(_2421_),
    .A2(_2422_),
    .ZN(_2423_));
 OAI22_X1 _3259_ (.A1(_0018_),
    .A2(_2352_),
    .B1(_2353_),
    .B2(_2265_),
    .ZN(_2424_));
 NOR2_X1 _3260_ (.A1(_2320_),
    .A2(_2348_),
    .ZN(_2425_));
 AOI21_X1 _3261_ (.A(_2425_),
    .B1(_2349_),
    .B2(_2351_),
    .ZN(_2426_));
 INV_X1 _3262_ (.A(_2345_),
    .ZN(_2427_));
 NOR2_X1 _3263_ (.A1(_2427_),
    .A2(_2347_),
    .ZN(_2428_));
 INV_X1 _3264_ (.A(net82),
    .ZN(_2429_));
 INV_X1 _3265_ (.A(net61),
    .ZN(_2430_));
 OR2_X1 _3266_ (.A1(_2430_),
    .A2(_2342_),
    .ZN(_2431_));
 INV_X1 _3267_ (.A(net85),
    .ZN(_2432_));
 NOR2_X1 _3268_ (.A1(_2326_),
    .A2(_2339_),
    .ZN(_2433_));
 NOR2_X1 _3269_ (.A1(_2330_),
    .A2(_2337_),
    .ZN(_2434_));
 AOI21_X1 _3270_ (.A(_2434_),
    .B1(_2338_),
    .B2(_2328_),
    .ZN(_2435_));
 NAND2_X1 _3271_ (.A1(\iir1.y[4] ),
    .A2(\iir1.y[2] ),
    .ZN(_2436_));
 AND2_X1 _3272_ (.A1(\iir1.y[4] ),
    .A2(_2279_),
    .ZN(_2437_));
 OAI21_X1 _3273_ (.A(_2334_),
    .B1(_2437_),
    .B2(_2331_),
    .ZN(_2438_));
 OAI21_X1 _3274_ (.A(_2438_),
    .B1(_2335_),
    .B2(_2336_),
    .ZN(_2439_));
 XOR2_X1 _3275_ (.A(\iir1.y[8] ),
    .B(\iir1.y[7] ),
    .Z(_2440_));
 XNOR2_X1 _3276_ (.A(\iir1.y[6] ),
    .B(_2440_),
    .ZN(_2441_));
 NAND2_X1 _3277_ (.A1(\iir1.y[7] ),
    .A2(\iir1.y[6] ),
    .ZN(_2442_));
 OAI21_X1 _3278_ (.A(\iir1.y[5] ),
    .B1(\iir1.y[6] ),
    .B2(\iir1.y[7] ),
    .ZN(_2443_));
 NAND2_X1 _3279_ (.A1(_2442_),
    .A2(_2443_),
    .ZN(_2444_));
 XNOR2_X1 _3280_ (.A(_2441_),
    .B(_2444_),
    .ZN(_2445_));
 XOR2_X1 _3281_ (.A(_1968_),
    .B(_2445_),
    .Z(_2446_));
 XNOR2_X1 _3282_ (.A(_2439_),
    .B(_2446_),
    .ZN(_2447_));
 XNOR2_X1 _3283_ (.A(_2436_),
    .B(_2447_),
    .ZN(_2448_));
 XOR2_X1 _3284_ (.A(_2435_),
    .B(_2448_),
    .Z(_2449_));
 XNOR2_X1 _3285_ (.A(_2433_),
    .B(_2449_),
    .ZN(_2450_));
 AND3_X1 _3286_ (.A1(_2285_),
    .A2(_2284_),
    .A3(_2340_),
    .ZN(_2451_));
 AOI21_X1 _3287_ (.A(_2451_),
    .B1(_2341_),
    .B2(_2323_),
    .ZN(_2452_));
 XNOR2_X1 _3288_ (.A(_2450_),
    .B(_2452_),
    .ZN(_2453_));
 XNOR2_X1 _3289_ (.A(_2432_),
    .B(_2453_),
    .ZN(_2454_));
 XOR2_X1 _3290_ (.A(_2431_),
    .B(_2454_),
    .Z(_2455_));
 XNOR2_X1 _3291_ (.A(_2429_),
    .B(_2455_),
    .ZN(_2456_));
 AND3_X1 _3292_ (.A1(\iir1.y2[5] ),
    .A2(_2288_),
    .A3(_2343_),
    .ZN(_2457_));
 AOI21_X1 _3293_ (.A(_2457_),
    .B1(_2344_),
    .B2(_0012_),
    .ZN(_2458_));
 XOR2_X1 _3294_ (.A(_2456_),
    .B(_2458_),
    .Z(_2459_));
 XNOR2_X1 _3295_ (.A(_2428_),
    .B(_2459_),
    .ZN(_2460_));
 XOR2_X1 _3296_ (.A(_2426_),
    .B(_2460_),
    .Z(_2461_));
 XNOR2_X1 _3297_ (.A(\iir2.x2[8] ),
    .B(_2461_),
    .ZN(_2462_));
 XOR2_X1 _3298_ (.A(_0018_),
    .B(_2462_),
    .Z(_2463_));
 XNOR2_X1 _3299_ (.A(_2424_),
    .B(_2463_),
    .ZN(_2464_));
 XNOR2_X1 _3300_ (.A(\iir2.x2[5] ),
    .B(\iir2.x2[6] ),
    .ZN(_2465_));
 XNOR2_X1 _3301_ (.A(_2464_),
    .B(_2465_),
    .ZN(_2466_));
 XNOR2_X1 _3302_ (.A(_2423_),
    .B(_2466_),
    .ZN(_2467_));
 NAND2_X1 _3303_ (.A1(\iir2.x2[4] ),
    .A2(\iir2.x2[5] ),
    .ZN(_2468_));
 XOR2_X1 _3304_ (.A(_0021_),
    .B(_2468_),
    .Z(_2469_));
 XNOR2_X1 _3305_ (.A(_2467_),
    .B(_2469_),
    .ZN(_2470_));
 XOR2_X1 _3306_ (.A(_2420_),
    .B(_2470_),
    .Z(_2471_));
 XNOR2_X1 _3307_ (.A(_2415_),
    .B(_2471_),
    .ZN(_2472_));
 XNOR2_X1 _3308_ (.A(_2414_),
    .B(_2472_),
    .ZN(_2473_));
 XOR2_X1 _3309_ (.A(_2412_),
    .B(_2473_),
    .Z(_2474_));
 NAND2_X1 _3310_ (.A1(z[5]),
    .A2(_2474_),
    .ZN(_2475_));
 AOI21_X1 _3311_ (.A(_2470_),
    .B1(_2419_),
    .B2(_2417_),
    .ZN(_2476_));
 NAND3_X1 _3312_ (.A1(_2417_),
    .A2(_2419_),
    .A3(_2470_),
    .ZN(_2477_));
 AOI21_X1 _3313_ (.A(_2476_),
    .B1(_2477_),
    .B2(_2415_),
    .ZN(_2478_));
 NOR2_X1 _3314_ (.A1(_0021_),
    .A2(_2468_),
    .ZN(_2479_));
 AOI21_X1 _3315_ (.A(_2466_),
    .B1(_2422_),
    .B2(_2421_),
    .ZN(_2480_));
 AOI21_X1 _3316_ (.A(_2480_),
    .B1(_2467_),
    .B2(_2469_),
    .ZN(_2481_));
 NAND2_X1 _3317_ (.A1(_2424_),
    .A2(_2463_),
    .ZN(_2482_));
 NOR2_X1 _3318_ (.A1(_2424_),
    .A2(_2463_),
    .ZN(_2483_));
 OAI21_X1 _3319_ (.A(_2482_),
    .B1(_2465_),
    .B2(_2483_),
    .ZN(_2484_));
 INV_X1 _3320_ (.A(_2461_),
    .ZN(_2485_));
 OAI22_X1 _3321_ (.A1(_0016_),
    .A2(_2485_),
    .B1(_2462_),
    .B2(_2319_),
    .ZN(_2486_));
 NAND2_X1 _3322_ (.A1(_2428_),
    .A2(_2459_),
    .ZN(_2487_));
 OAI21_X1 _3323_ (.A(_2487_),
    .B1(_2460_),
    .B2(_2426_),
    .ZN(_2488_));
 NOR2_X1 _3324_ (.A1(_2456_),
    .A2(_2458_),
    .ZN(_2489_));
 OR2_X1 _3325_ (.A1(_2432_),
    .A2(_2453_),
    .ZN(_2490_));
 INV_X1 _3326_ (.A(net70),
    .ZN(_2491_));
 NOR2_X1 _3327_ (.A1(_2435_),
    .A2(_2448_),
    .ZN(_2492_));
 NAND2_X1 _3328_ (.A1(_2439_),
    .A2(_2446_),
    .ZN(_2493_));
 OAI21_X1 _3329_ (.A(_2493_),
    .B1(_2447_),
    .B2(_2436_),
    .ZN(_2494_));
 AND2_X1 _3330_ (.A1(\iir1.y[5] ),
    .A2(\iir1.y[3] ),
    .ZN(_2495_));
 AOI21_X1 _3331_ (.A(_2441_),
    .B1(_2443_),
    .B2(_2442_),
    .ZN(_2496_));
 AOI21_X1 _3332_ (.A(_2496_),
    .B1(_2445_),
    .B2(_1968_),
    .ZN(_2497_));
 AND2_X1 _3333_ (.A1(\iir1.y[8] ),
    .A2(\iir1.y[7] ),
    .ZN(_2498_));
 AOI21_X1 _3334_ (.A(_2498_),
    .B1(_2440_),
    .B2(\iir1.y[6] ),
    .ZN(_2499_));
 XOR2_X1 _3335_ (.A(\iir1.y[9] ),
    .B(\iir1.y[8] ),
    .Z(_2500_));
 XNOR2_X1 _3336_ (.A(\iir1.y[7] ),
    .B(_2500_),
    .ZN(_2501_));
 XOR2_X1 _3337_ (.A(_2499_),
    .B(_2501_),
    .Z(_2502_));
 XNOR2_X1 _3338_ (.A(\iir1.y[6] ),
    .B(\iir1.y[4] ),
    .ZN(_2503_));
 INV_X1 _3339_ (.A(_2503_),
    .ZN(_2504_));
 XNOR2_X1 _3340_ (.A(_2502_),
    .B(_2504_),
    .ZN(_2505_));
 XOR2_X1 _3341_ (.A(_2497_),
    .B(_2505_),
    .Z(_2506_));
 XOR2_X1 _3342_ (.A(_2495_),
    .B(_2506_),
    .Z(_2507_));
 XOR2_X1 _3343_ (.A(_2494_),
    .B(_2507_),
    .Z(_2508_));
 XNOR2_X1 _3344_ (.A(_2492_),
    .B(_2508_),
    .ZN(_2509_));
 NAND2_X1 _3345_ (.A1(_2433_),
    .A2(_2449_),
    .ZN(_2510_));
 OAI21_X1 _3346_ (.A(_2510_),
    .B1(_2450_),
    .B2(_2452_),
    .ZN(_2511_));
 XOR2_X1 _3347_ (.A(_2509_),
    .B(_2511_),
    .Z(_2512_));
 XNOR2_X1 _3348_ (.A(_2491_),
    .B(_2512_),
    .ZN(_2513_));
 XOR2_X1 _3349_ (.A(_2490_),
    .B(_2513_),
    .Z(_2514_));
 XNOR2_X1 _3350_ (.A(_0009_),
    .B(_2514_),
    .ZN(_2515_));
 NOR2_X1 _3351_ (.A1(_2431_),
    .A2(_2454_),
    .ZN(_2516_));
 AOI21_X1 _3352_ (.A(_2516_),
    .B1(_2455_),
    .B2(_0011_),
    .ZN(_2517_));
 XNOR2_X1 _3353_ (.A(_2515_),
    .B(_2517_),
    .ZN(_2518_));
 XNOR2_X1 _3354_ (.A(_2489_),
    .B(_2518_),
    .ZN(_2519_));
 XNOR2_X1 _3355_ (.A(_2488_),
    .B(_2519_),
    .ZN(_2520_));
 XNOR2_X1 _3356_ (.A(_0016_),
    .B(\iir2.x2[9] ),
    .ZN(_2521_));
 XNOR2_X1 _3357_ (.A(_2520_),
    .B(_2521_),
    .ZN(_2522_));
 XNOR2_X1 _3358_ (.A(_2486_),
    .B(_2522_),
    .ZN(_2523_));
 XNOR2_X1 _3359_ (.A(\iir2.x2[7] ),
    .B(\iir2.x2[6] ),
    .ZN(_2524_));
 XOR2_X1 _3360_ (.A(_2523_),
    .B(_2524_),
    .Z(_2525_));
 XNOR2_X1 _3361_ (.A(_2484_),
    .B(_2525_),
    .ZN(_2526_));
 NAND2_X1 _3362_ (.A1(\iir2.x2[5] ),
    .A2(\iir2.x2[6] ),
    .ZN(_2527_));
 XNOR2_X1 _3363_ (.A(_0019_),
    .B(_2527_),
    .ZN(_2528_));
 XOR2_X1 _3364_ (.A(_2526_),
    .B(_2528_),
    .Z(_2529_));
 XNOR2_X1 _3365_ (.A(_2481_),
    .B(_2529_),
    .ZN(_2530_));
 XNOR2_X1 _3366_ (.A(_2479_),
    .B(_2530_),
    .ZN(_2531_));
 XNOR2_X1 _3367_ (.A(_2478_),
    .B(_2531_),
    .ZN(_2532_));
 NAND2_X1 _3368_ (.A1(_2414_),
    .A2(_2472_),
    .ZN(_2533_));
 OAI21_X1 _3369_ (.A(_2533_),
    .B1(_2473_),
    .B2(_2412_),
    .ZN(_2534_));
 XNOR2_X1 _3370_ (.A(_2532_),
    .B(_2534_),
    .ZN(_2535_));
 XNOR2_X1 _3371_ (.A(z[6]),
    .B(_2535_),
    .ZN(_2536_));
 NOR2_X1 _3372_ (.A1(_2475_),
    .A2(_2536_),
    .ZN(_2537_));
 NAND2_X1 _3373_ (.A1(z[6]),
    .A2(_2535_),
    .ZN(_2538_));
 NOR3_X1 _3374_ (.A1(_2412_),
    .A2(_2473_),
    .A3(_2532_),
    .ZN(_2539_));
 OR2_X1 _3375_ (.A1(_2478_),
    .A2(_2531_),
    .ZN(_2540_));
 OAI21_X1 _3376_ (.A(_2540_),
    .B1(_2532_),
    .B2(_2533_),
    .ZN(_2541_));
 OR2_X1 _3377_ (.A1(_2539_),
    .A2(_2541_),
    .ZN(_2542_));
 INV_X1 _3378_ (.A(_2529_),
    .ZN(_2543_));
 NOR2_X1 _3379_ (.A1(_2481_),
    .A2(_2543_),
    .ZN(_2544_));
 AOI21_X1 _3380_ (.A(_2544_),
    .B1(_2530_),
    .B2(_2479_),
    .ZN(_2545_));
 NOR2_X1 _3381_ (.A1(_0019_),
    .A2(_2527_),
    .ZN(_2546_));
 NOR2_X1 _3382_ (.A1(_2526_),
    .A2(_2528_),
    .ZN(_2547_));
 AOI21_X1 _3383_ (.A(_2547_),
    .B1(_2525_),
    .B2(_2484_),
    .ZN(_2548_));
 NAND2_X1 _3384_ (.A1(\iir2.x2[7] ),
    .A2(\iir2.x2[6] ),
    .ZN(_2549_));
 XOR2_X1 _3385_ (.A(_0017_),
    .B(_2549_),
    .Z(_2550_));
 NOR2_X1 _3386_ (.A1(_2523_),
    .A2(_2524_),
    .ZN(_2551_));
 AOI21_X1 _3387_ (.A(_2551_),
    .B1(_2522_),
    .B2(_2486_),
    .ZN(_2552_));
 XOR2_X1 _3388_ (.A(\iir2.x2[8] ),
    .B(\iir2.x2[7] ),
    .Z(_2553_));
 INV_X1 _3389_ (.A(\iir2.x2[10] ),
    .ZN(_2554_));
 NOR3_X1 _3390_ (.A1(_2456_),
    .A2(_2458_),
    .A3(_2518_),
    .ZN(_2555_));
 AOI21_X1 _3391_ (.A(_2555_),
    .B1(_2519_),
    .B2(_2488_),
    .ZN(_2556_));
 NOR2_X1 _3392_ (.A1(_2515_),
    .A2(_2517_),
    .ZN(_2557_));
 NOR2_X1 _3393_ (.A1(_2490_),
    .A2(_2513_),
    .ZN(_2558_));
 AOI21_X1 _3394_ (.A(_2558_),
    .B1(_2514_),
    .B2(_0009_),
    .ZN(_2559_));
 NOR2_X1 _3395_ (.A1(_0008_),
    .A2(_2512_),
    .ZN(_2560_));
 INV_X1 _3396_ (.A(net87),
    .ZN(_2561_));
 NAND2_X1 _3397_ (.A1(_2492_),
    .A2(_2508_),
    .ZN(_2562_));
 OR2_X1 _3398_ (.A1(_2450_),
    .A2(_2509_),
    .ZN(_2563_));
 OAI221_X1 _3399_ (.A(_2562_),
    .B1(_2509_),
    .B2(_2510_),
    .C1(_2563_),
    .C2(_2452_),
    .ZN(_2564_));
 NAND2_X1 _3400_ (.A1(_2494_),
    .A2(_2507_),
    .ZN(_2565_));
 NOR2_X1 _3401_ (.A1(_2497_),
    .A2(_2505_),
    .ZN(_2566_));
 AOI21_X1 _3402_ (.A(_2566_),
    .B1(_2506_),
    .B2(_2495_),
    .ZN(_2567_));
 AND2_X1 _3403_ (.A1(\iir1.y[6] ),
    .A2(\iir1.y[4] ),
    .ZN(_2568_));
 NOR2_X1 _3404_ (.A1(_2499_),
    .A2(_2501_),
    .ZN(_2569_));
 AOI21_X1 _3405_ (.A(_2569_),
    .B1(_2502_),
    .B2(_2504_),
    .ZN(_2570_));
 XNOR2_X1 _3406_ (.A(\iir1.y[7] ),
    .B(\iir1.y[5] ),
    .ZN(_2571_));
 XNOR2_X1 _3407_ (.A(\iir1.y[9] ),
    .B(\iir1.y[10] ),
    .ZN(_2572_));
 XOR2_X1 _3408_ (.A(\iir1.y[8] ),
    .B(_2572_),
    .Z(_2573_));
 AND2_X1 _3409_ (.A1(\iir1.y[9] ),
    .A2(\iir1.y[8] ),
    .ZN(_2574_));
 AOI21_X1 _3410_ (.A(_2574_),
    .B1(_2500_),
    .B2(\iir1.y[7] ),
    .ZN(_2575_));
 XNOR2_X1 _3411_ (.A(_2573_),
    .B(_2575_),
    .ZN(_2576_));
 XNOR2_X1 _3412_ (.A(_2571_),
    .B(_2576_),
    .ZN(_2577_));
 XOR2_X1 _3413_ (.A(_2570_),
    .B(_2577_),
    .Z(_2578_));
 XOR2_X1 _3414_ (.A(_2568_),
    .B(_2578_),
    .Z(_2579_));
 XNOR2_X1 _3415_ (.A(_2567_),
    .B(_2579_),
    .ZN(_2580_));
 XOR2_X1 _3416_ (.A(_2565_),
    .B(_2580_),
    .Z(_2581_));
 INV_X1 _3417_ (.A(_2581_),
    .ZN(_2582_));
 XNOR2_X1 _3418_ (.A(_2564_),
    .B(_2582_),
    .ZN(_2583_));
 XNOR2_X1 _3419_ (.A(_2561_),
    .B(_2583_),
    .ZN(_2584_));
 XNOR2_X1 _3420_ (.A(_2560_),
    .B(_2584_),
    .ZN(_2585_));
 XNOR2_X1 _3421_ (.A(_0003_),
    .B(_2585_),
    .ZN(_2586_));
 XOR2_X1 _3422_ (.A(_2559_),
    .B(_2586_),
    .Z(_2587_));
 XOR2_X1 _3423_ (.A(_2557_),
    .B(_2587_),
    .Z(_2588_));
 XNOR2_X1 _3424_ (.A(_2556_),
    .B(_2588_),
    .ZN(_2589_));
 XNOR2_X1 _3425_ (.A(_2554_),
    .B(_2589_),
    .ZN(_2590_));
 XNOR2_X1 _3426_ (.A(\iir2.x2[9] ),
    .B(_2590_),
    .ZN(_2591_));
 NOR2_X1 _3427_ (.A1(\iir2.x2[9] ),
    .A2(\iir2.x2[8] ),
    .ZN(_2592_));
 NOR2_X1 _3428_ (.A1(_2520_),
    .A2(_2592_),
    .ZN(_2593_));
 AOI21_X1 _3429_ (.A(_2593_),
    .B1(\iir2.x2[8] ),
    .B2(\iir2.x2[9] ),
    .ZN(_2594_));
 XOR2_X1 _3430_ (.A(_2591_),
    .B(_2594_),
    .Z(_2595_));
 XNOR2_X1 _3431_ (.A(_2553_),
    .B(_2595_),
    .ZN(_2596_));
 XOR2_X1 _3432_ (.A(_2552_),
    .B(_2596_),
    .Z(_2597_));
 XNOR2_X1 _3433_ (.A(_2550_),
    .B(_2597_),
    .ZN(_2598_));
 XOR2_X1 _3434_ (.A(_2548_),
    .B(_2598_),
    .Z(_2599_));
 XNOR2_X1 _3435_ (.A(_2546_),
    .B(_2599_),
    .ZN(_2600_));
 XOR2_X1 _3436_ (.A(_2545_),
    .B(_2600_),
    .Z(_2601_));
 XOR2_X1 _3437_ (.A(_2542_),
    .B(_2601_),
    .Z(_2602_));
 XNOR2_X1 _3438_ (.A(z[7]),
    .B(_2602_),
    .ZN(_2603_));
 XOR2_X1 _3439_ (.A(_2538_),
    .B(_2603_),
    .Z(_2604_));
 XNOR2_X1 _3440_ (.A(_2537_),
    .B(_2604_),
    .ZN(_2605_));
 NOR2_X1 _3441_ (.A1(_1330_),
    .A2(_2605_),
    .ZN(_2606_));
 AOI21_X1 _3442_ (.A(_2606_),
    .B1(_2604_),
    .B2(_2537_),
    .ZN(_2607_));
 NAND2_X1 _3443_ (.A1(z[1]),
    .A2(z[0]),
    .ZN(_2608_));
 XOR2_X1 _3444_ (.A(z[2]),
    .B(z[1]),
    .Z(_2609_));
 XNOR2_X1 _3445_ (.A(_2608_),
    .B(_2609_),
    .ZN(_2610_));
 NOR2_X1 _3446_ (.A1(_2538_),
    .A2(_2603_),
    .ZN(_2611_));
 AND2_X1 _3447_ (.A1(z[7]),
    .A2(_2602_),
    .ZN(_2612_));
 INV_X1 _3448_ (.A(net74),
    .ZN(_2613_));
 NOR2_X1 _3449_ (.A1(_2545_),
    .A2(_2600_),
    .ZN(_2614_));
 AOI21_X1 _3450_ (.A(_2614_),
    .B1(_2601_),
    .B2(_2542_),
    .ZN(_2615_));
 NOR2_X1 _3451_ (.A1(_2548_),
    .A2(_2598_),
    .ZN(_2616_));
 AOI21_X1 _3452_ (.A(_2616_),
    .B1(_2599_),
    .B2(_2546_),
    .ZN(_2617_));
 NOR2_X1 _3453_ (.A1(_0017_),
    .A2(_2549_),
    .ZN(_2618_));
 NOR2_X1 _3454_ (.A1(_2552_),
    .A2(_2596_),
    .ZN(_2619_));
 AOI21_X1 _3455_ (.A(_2619_),
    .B1(_2597_),
    .B2(_2550_),
    .ZN(_2620_));
 NAND2_X1 _3456_ (.A1(\iir2.x2[8] ),
    .A2(\iir2.x2[7] ),
    .ZN(_2621_));
 XNOR2_X1 _3457_ (.A(_2316_),
    .B(_2621_),
    .ZN(_2622_));
 NOR2_X1 _3458_ (.A1(_2591_),
    .A2(_2594_),
    .ZN(_2623_));
 AOI21_X1 _3459_ (.A(_2623_),
    .B1(_2595_),
    .B2(_2553_),
    .ZN(_2624_));
 XNOR2_X1 _3460_ (.A(\iir2.x2[9] ),
    .B(\iir2.x2[8] ),
    .ZN(_2625_));
 INV_X1 _3461_ (.A(_0031_),
    .ZN(_2626_));
 AOI22_X1 _3462_ (.A1(_2626_),
    .A2(_2589_),
    .B1(_2590_),
    .B2(\iir2.x2[9] ),
    .ZN(_2627_));
 NAND3_X1 _3463_ (.A1(_2488_),
    .A2(_2519_),
    .A3(_2588_),
    .ZN(_2628_));
 AND2_X1 _3464_ (.A1(_2557_),
    .A2(_2587_),
    .ZN(_2629_));
 AOI21_X1 _3465_ (.A(_2629_),
    .B1(_2588_),
    .B2(_2555_),
    .ZN(_2630_));
 AND2_X1 _3466_ (.A1(_2628_),
    .A2(_2630_),
    .ZN(_2631_));
 NOR2_X1 _3467_ (.A1(_2559_),
    .A2(_2586_),
    .ZN(_2632_));
 INV_X1 _3468_ (.A(_2632_),
    .ZN(_2633_));
 NOR3_X1 _3469_ (.A1(_0008_),
    .A2(_2512_),
    .A3(_2584_),
    .ZN(_2634_));
 AOI21_X1 _3470_ (.A(_2634_),
    .B1(_2585_),
    .B2(_0003_),
    .ZN(_2635_));
 NOR2_X1 _3471_ (.A1(_0030_),
    .A2(_2583_),
    .ZN(_2636_));
 AND3_X1 _3472_ (.A1(_2494_),
    .A2(_2507_),
    .A3(_2580_),
    .ZN(_2637_));
 AOI21_X1 _3473_ (.A(_2637_),
    .B1(_2582_),
    .B2(_2564_),
    .ZN(_2638_));
 AND2_X1 _3474_ (.A1(_2495_),
    .A2(_2506_),
    .ZN(_2639_));
 OAI21_X1 _3475_ (.A(_2579_),
    .B1(_2639_),
    .B2(_2566_),
    .ZN(_2640_));
 NOR2_X1 _3476_ (.A1(_2570_),
    .A2(_2577_),
    .ZN(_2641_));
 AOI21_X1 _3477_ (.A(_2641_),
    .B1(_2578_),
    .B2(_2568_),
    .ZN(_2642_));
 NAND2_X1 _3478_ (.A1(\iir1.y[7] ),
    .A2(\iir1.y[5] ),
    .ZN(_2643_));
 OR2_X1 _3479_ (.A1(_2573_),
    .A2(_2575_),
    .ZN(_2644_));
 OAI21_X1 _3480_ (.A(_2644_),
    .B1(_2576_),
    .B2(_2571_),
    .ZN(_2645_));
 XOR2_X1 _3481_ (.A(\iir1.y[8] ),
    .B(\iir1.y[6] ),
    .Z(_2646_));
 AND2_X1 _3482_ (.A1(\iir1.y[8] ),
    .A2(\iir1.y[10] ),
    .ZN(_2647_));
 OR2_X1 _3483_ (.A1(\iir1.y[9] ),
    .A2(_2647_),
    .ZN(_2648_));
 OAI21_X1 _3484_ (.A(\iir1.y[9] ),
    .B1(\iir1.y[8] ),
    .B2(\iir1.y[10] ),
    .ZN(_2649_));
 NAND2_X1 _3485_ (.A1(_2648_),
    .A2(_2649_),
    .ZN(_2650_));
 XNOR2_X1 _3486_ (.A(_2646_),
    .B(_2650_),
    .ZN(_2651_));
 XNOR2_X1 _3487_ (.A(_2645_),
    .B(_2651_),
    .ZN(_2652_));
 XOR2_X1 _3488_ (.A(_2643_),
    .B(_2652_),
    .Z(_2653_));
 XNOR2_X1 _3489_ (.A(_2642_),
    .B(_2653_),
    .ZN(_2654_));
 XOR2_X1 _3490_ (.A(_2640_),
    .B(_2654_),
    .Z(_2655_));
 INV_X1 _3491_ (.A(_2655_),
    .ZN(_2656_));
 XNOR2_X1 _3492_ (.A(_2638_),
    .B(_2656_),
    .ZN(_2657_));
 XNOR2_X1 _3493_ (.A(\iir1.y2[10] ),
    .B(_2657_),
    .ZN(_2658_));
 XNOR2_X1 _3494_ (.A(_2636_),
    .B(_2658_),
    .ZN(_2659_));
 XNOR2_X1 _3495_ (.A(_2432_),
    .B(_2659_),
    .ZN(_2660_));
 XNOR2_X1 _3496_ (.A(_2635_),
    .B(_2660_),
    .ZN(_2661_));
 XNOR2_X1 _3497_ (.A(_2633_),
    .B(_2661_),
    .ZN(_2662_));
 XNOR2_X1 _3498_ (.A(_2631_),
    .B(_2662_),
    .ZN(_2663_));
 XNOR2_X1 _3499_ (.A(_2627_),
    .B(_2663_),
    .ZN(_2664_));
 XNOR2_X1 _3500_ (.A(_2625_),
    .B(_2664_),
    .ZN(_2665_));
 XOR2_X1 _3501_ (.A(_2624_),
    .B(_2665_),
    .Z(_2666_));
 XNOR2_X1 _3502_ (.A(_2622_),
    .B(_2666_),
    .ZN(_2667_));
 XOR2_X1 _3503_ (.A(_2620_),
    .B(_2667_),
    .Z(_2668_));
 XNOR2_X1 _3504_ (.A(_2618_),
    .B(_2668_),
    .ZN(_2669_));
 XOR2_X1 _3505_ (.A(_2617_),
    .B(_2669_),
    .Z(_2670_));
 XNOR2_X1 _3506_ (.A(_2615_),
    .B(_2670_),
    .ZN(_2671_));
 XNOR2_X1 _3507_ (.A(_2613_),
    .B(_2671_),
    .ZN(_2672_));
 XOR2_X1 _3508_ (.A(_2612_),
    .B(_2672_),
    .Z(_2673_));
 XOR2_X1 _3509_ (.A(_2611_),
    .B(_2673_),
    .Z(_2674_));
 XNOR2_X1 _3510_ (.A(_2610_),
    .B(_2674_),
    .ZN(_2675_));
 OR2_X1 _3511_ (.A1(_2607_),
    .A2(_2675_),
    .ZN(_2676_));
 INV_X1 _3512_ (.A(_2676_),
    .ZN(_2677_));
 NOR2_X1 _3513_ (.A1(z[2]),
    .A2(_2608_),
    .ZN(_2678_));
 AND2_X1 _3514_ (.A1(_2611_),
    .A2(_2673_),
    .ZN(_2679_));
 AOI21_X1 _3515_ (.A(_2679_),
    .B1(_2674_),
    .B2(_2610_),
    .ZN(_2680_));
 NAND2_X1 _3516_ (.A1(z[2]),
    .A2(z[1]),
    .ZN(_2681_));
 XOR2_X1 _3517_ (.A(z[3]),
    .B(z[2]),
    .Z(_2682_));
 XNOR2_X1 _3518_ (.A(_2681_),
    .B(_2682_),
    .ZN(_2683_));
 NAND2_X1 _3519_ (.A1(_2612_),
    .A2(_2672_),
    .ZN(_2684_));
 NAND2_X1 _3520_ (.A1(z[8]),
    .A2(_2671_),
    .ZN(_2685_));
 NOR2_X1 _3521_ (.A1(_2617_),
    .A2(_2669_),
    .ZN(_2686_));
 AOI21_X1 _3522_ (.A(_2686_),
    .B1(_2670_),
    .B2(_2614_),
    .ZN(_2687_));
 NAND3_X1 _3523_ (.A1(_2542_),
    .A2(_2601_),
    .A3(_2670_),
    .ZN(_2688_));
 NOR2_X1 _3524_ (.A1(_2620_),
    .A2(_2667_),
    .ZN(_2689_));
 AOI21_X1 _3525_ (.A(_2689_),
    .B1(_2668_),
    .B2(_2618_),
    .ZN(_2690_));
 NOR2_X1 _3526_ (.A1(_0020_),
    .A2(_2621_),
    .ZN(_2691_));
 NOR2_X1 _3527_ (.A1(_2624_),
    .A2(_2665_),
    .ZN(_2692_));
 AOI21_X1 _3528_ (.A(_2692_),
    .B1(_2666_),
    .B2(_2622_),
    .ZN(_2693_));
 NAND2_X1 _3529_ (.A1(\iir2.x2[9] ),
    .A2(\iir2.x2[8] ),
    .ZN(_2694_));
 XOR2_X1 _3530_ (.A(_0018_),
    .B(_2694_),
    .Z(_2695_));
 OR2_X1 _3531_ (.A1(_2627_),
    .A2(_2663_),
    .ZN(_2696_));
 OAI21_X1 _3532_ (.A(_2696_),
    .B1(_2664_),
    .B2(_2625_),
    .ZN(_2697_));
 XOR2_X1 _3533_ (.A(\iir2.x2[10] ),
    .B(\iir2.x2[9] ),
    .Z(_2698_));
 INV_X1 _3534_ (.A(_2698_),
    .ZN(_2699_));
 NOR2_X1 _3535_ (.A1(_2633_),
    .A2(_2661_),
    .ZN(_2700_));
 INV_X1 _3536_ (.A(_2700_),
    .ZN(_2701_));
 OAI21_X1 _3537_ (.A(_2701_),
    .B1(_2662_),
    .B2(_2631_),
    .ZN(_2702_));
 NOR2_X1 _3538_ (.A1(_2635_),
    .A2(_2660_),
    .ZN(_2703_));
 INV_X1 _3539_ (.A(\iir1.y2[10] ),
    .ZN(_2704_));
 NOR2_X1 _3540_ (.A1(_2704_),
    .A2(_2657_),
    .ZN(_2705_));
 OR4_X1 _3541_ (.A1(_2452_),
    .A2(_2563_),
    .A3(_2581_),
    .A4(_2655_),
    .ZN(_2706_));
 INV_X1 _3542_ (.A(_2654_),
    .ZN(_2707_));
 NOR2_X1 _3543_ (.A1(_2640_),
    .A2(_2707_),
    .ZN(_2708_));
 NOR2_X1 _3544_ (.A1(_2581_),
    .A2(_2655_),
    .ZN(_2709_));
 OAI21_X1 _3545_ (.A(_2562_),
    .B1(_2509_),
    .B2(_2510_),
    .ZN(_2710_));
 AOI221_X1 _3546_ (.A(_2708_),
    .B1(_2656_),
    .B2(_2637_),
    .C1(_2709_),
    .C2(_2710_),
    .ZN(_2711_));
 NAND2_X1 _3547_ (.A1(_2706_),
    .A2(_2711_),
    .ZN(_2712_));
 INV_X1 _3548_ (.A(_2653_),
    .ZN(_2713_));
 NOR2_X1 _3549_ (.A1(_2642_),
    .A2(_2713_),
    .ZN(_2714_));
 NOR2_X1 _3550_ (.A1(_2643_),
    .A2(_2652_),
    .ZN(_2715_));
 AOI21_X1 _3551_ (.A(_2715_),
    .B1(_2651_),
    .B2(_2645_),
    .ZN(_2716_));
 NAND2_X1 _3552_ (.A1(\iir1.y[8] ),
    .A2(\iir1.y[6] ),
    .ZN(_2717_));
 XOR2_X1 _3553_ (.A(\iir1.y[9] ),
    .B(\iir1.y[7] ),
    .Z(_2718_));
 NAND3_X1 _3554_ (.A1(_2646_),
    .A2(_2648_),
    .A3(_2649_),
    .ZN(_2719_));
 NAND2_X1 _3555_ (.A1(\iir1.y[9] ),
    .A2(\iir1.y[10] ),
    .ZN(_2720_));
 NAND2_X1 _3556_ (.A1(\iir1.y[8] ),
    .A2(\iir1.y[10] ),
    .ZN(_2721_));
 NAND2_X1 _3557_ (.A1(_2720_),
    .A2(_2721_),
    .ZN(_2722_));
 NOR2_X1 _3558_ (.A1(_2574_),
    .A2(_2722_),
    .ZN(_2723_));
 OAI21_X1 _3559_ (.A(_2719_),
    .B1(_2723_),
    .B2(_0000_),
    .ZN(_2724_));
 XOR2_X1 _3560_ (.A(_2718_),
    .B(_2724_),
    .Z(_2725_));
 XNOR2_X1 _3561_ (.A(_2717_),
    .B(_2725_),
    .ZN(_2726_));
 XNOR2_X1 _3562_ (.A(_2716_),
    .B(_2726_),
    .ZN(_2727_));
 XOR2_X1 _3563_ (.A(_2714_),
    .B(_2727_),
    .Z(_2728_));
 XOR2_X1 _3564_ (.A(_2712_),
    .B(_2728_),
    .Z(_2729_));
 XOR2_X1 _3565_ (.A(_2705_),
    .B(_2729_),
    .Z(_2730_));
 XOR2_X1 _3566_ (.A(_0008_),
    .B(_2730_),
    .Z(_2731_));
 NOR3_X1 _3567_ (.A1(_0030_),
    .A2(_2583_),
    .A3(_2658_),
    .ZN(_2732_));
 AOI21_X1 _3568_ (.A(_2732_),
    .B1(_2659_),
    .B2(_0001_),
    .ZN(_2733_));
 XNOR2_X1 _3569_ (.A(_2731_),
    .B(_2733_),
    .ZN(_2734_));
 XNOR2_X1 _3570_ (.A(_2703_),
    .B(_2734_),
    .ZN(_2735_));
 XNOR2_X1 _3571_ (.A(_2702_),
    .B(_2735_),
    .ZN(_2736_));
 XNOR2_X1 _3572_ (.A(_0031_),
    .B(_2736_),
    .ZN(_2737_));
 XNOR2_X1 _3573_ (.A(_2699_),
    .B(_2737_),
    .ZN(_2738_));
 XOR2_X1 _3574_ (.A(_2697_),
    .B(_2738_),
    .Z(_2739_));
 XNOR2_X1 _3575_ (.A(_2695_),
    .B(_2739_),
    .ZN(_2740_));
 XOR2_X1 _3576_ (.A(_2693_),
    .B(_2740_),
    .Z(_2741_));
 XNOR2_X1 _3577_ (.A(_2691_),
    .B(_2741_),
    .ZN(_2742_));
 XOR2_X1 _3578_ (.A(_2690_),
    .B(_2742_),
    .Z(_2743_));
 INV_X1 _3579_ (.A(_2743_),
    .ZN(_2744_));
 NAND3_X1 _3580_ (.A1(_2687_),
    .A2(_2688_),
    .A3(_2744_),
    .ZN(_2745_));
 AND3_X1 _3581_ (.A1(_2542_),
    .A2(_2601_),
    .A3(_2670_),
    .ZN(_2746_));
 OR2_X1 _3582_ (.A1(_2617_),
    .A2(_2669_),
    .ZN(_2747_));
 AND2_X1 _3583_ (.A1(_2617_),
    .A2(_2669_),
    .ZN(_2748_));
 OR2_X1 _3584_ (.A1(_2545_),
    .A2(_2600_),
    .ZN(_2749_));
 OAI21_X1 _3585_ (.A(_2747_),
    .B1(_2748_),
    .B2(_2749_),
    .ZN(_2750_));
 OAI21_X1 _3586_ (.A(_2743_),
    .B1(_2746_),
    .B2(_2750_),
    .ZN(_2751_));
 AOI21_X1 _3587_ (.A(z[9]),
    .B1(_2745_),
    .B2(_2751_),
    .ZN(_2752_));
 INV_X1 _3588_ (.A(net63),
    .ZN(_2753_));
 NOR3_X1 _3589_ (.A1(_2750_),
    .A2(_2746_),
    .A3(_2743_),
    .ZN(_2754_));
 AOI21_X1 _3590_ (.A(_2744_),
    .B1(_2688_),
    .B2(_2687_),
    .ZN(_2755_));
 NOR3_X1 _3591_ (.A1(_2753_),
    .A2(_2754_),
    .A3(_2755_),
    .ZN(_2756_));
 NOR3_X1 _3592_ (.A1(_2685_),
    .A2(_2752_),
    .A3(_2756_),
    .ZN(_2757_));
 AND2_X1 _3593_ (.A1(z[8]),
    .A2(_2671_),
    .ZN(_2758_));
 OAI21_X1 _3594_ (.A(_2753_),
    .B1(_2754_),
    .B2(_2755_),
    .ZN(_2759_));
 NAND3_X1 _3595_ (.A1(z[9]),
    .A2(_2745_),
    .A3(_2751_),
    .ZN(_2760_));
 AOI21_X1 _3596_ (.A(_2758_),
    .B1(_2759_),
    .B2(_2760_),
    .ZN(_2761_));
 OR3_X1 _3597_ (.A1(_2684_),
    .A2(_2757_),
    .A3(_2761_),
    .ZN(_2762_));
 OAI21_X1 _3598_ (.A(_2684_),
    .B1(_2757_),
    .B2(_2761_),
    .ZN(_2763_));
 AOI21_X1 _3599_ (.A(_2683_),
    .B1(_2762_),
    .B2(_2763_),
    .ZN(_2764_));
 INV_X1 _3600_ (.A(_2683_),
    .ZN(_2765_));
 NOR3_X1 _3601_ (.A1(_2684_),
    .A2(_2757_),
    .A3(_2761_),
    .ZN(_2766_));
 NAND3_X1 _3602_ (.A1(_2758_),
    .A2(_2759_),
    .A3(_2760_),
    .ZN(_2767_));
 OAI21_X1 _3603_ (.A(_2685_),
    .B1(_2752_),
    .B2(_2756_),
    .ZN(_2768_));
 AOI22_X1 _3604_ (.A1(_2612_),
    .A2(_2672_),
    .B1(_2767_),
    .B2(_2768_),
    .ZN(_2769_));
 NOR3_X1 _3605_ (.A1(_2765_),
    .A2(_2766_),
    .A3(_2769_),
    .ZN(_2770_));
 OR3_X1 _3606_ (.A1(_2680_),
    .A2(_2764_),
    .A3(_2770_),
    .ZN(_2771_));
 OAI21_X1 _3607_ (.A(_2680_),
    .B1(_2764_),
    .B2(_2770_),
    .ZN(_2772_));
 NAND3_X1 _3608_ (.A1(_2678_),
    .A2(_2771_),
    .A3(_2772_),
    .ZN(_2773_));
 NOR3_X1 _3609_ (.A1(_2680_),
    .A2(_2764_),
    .A3(_2770_),
    .ZN(_2774_));
 OAI21_X1 _3610_ (.A(_2765_),
    .B1(_2766_),
    .B2(_2769_),
    .ZN(_2775_));
 NAND3_X1 _3611_ (.A1(_2683_),
    .A2(_2762_),
    .A3(_2763_),
    .ZN(_2776_));
 AOI221_X1 _3612_ (.A(_2679_),
    .B1(_2775_),
    .B2(_2776_),
    .C1(_2674_),
    .C2(_2610_),
    .ZN(_2777_));
 OAI22_X1 _3613_ (.A1(z[2]),
    .A2(_2608_),
    .B1(_2774_),
    .B2(_2777_),
    .ZN(_2778_));
 NAND3_X1 _3614_ (.A1(_2677_),
    .A2(_2773_),
    .A3(_2778_),
    .ZN(_2779_));
 NAND2_X1 _3615_ (.A1(_2771_),
    .A2(_2773_),
    .ZN(_2780_));
 OR2_X1 _3616_ (.A1(z[3]),
    .A2(_2681_),
    .ZN(_2781_));
 NAND2_X1 _3617_ (.A1(_2762_),
    .A2(_2776_),
    .ZN(_2782_));
 NAND2_X1 _3618_ (.A1(z[3]),
    .A2(z[2]),
    .ZN(_2783_));
 XOR2_X1 _3619_ (.A(z[4]),
    .B(z[3]),
    .Z(_2784_));
 XNOR2_X1 _3620_ (.A(_2783_),
    .B(_2784_),
    .ZN(_2785_));
 INV_X1 _3621_ (.A(net75),
    .ZN(_2786_));
 NOR2_X1 _3622_ (.A1(_2693_),
    .A2(_2740_),
    .ZN(_2787_));
 AOI21_X1 _3623_ (.A(_2787_),
    .B1(_2741_),
    .B2(_2691_),
    .ZN(_2788_));
 OR2_X1 _3624_ (.A1(_0018_),
    .A2(_2694_),
    .ZN(_2789_));
 AND2_X1 _3625_ (.A1(_2697_),
    .A2(_2738_),
    .ZN(_2790_));
 AOI21_X1 _3626_ (.A(_2790_),
    .B1(_2739_),
    .B2(_2695_),
    .ZN(_2791_));
 NAND2_X1 _3627_ (.A1(\iir2.x2[10] ),
    .A2(\iir2.x2[9] ),
    .ZN(_2792_));
 XOR2_X1 _3628_ (.A(_0016_),
    .B(_2792_),
    .Z(_2793_));
 NAND2_X1 _3629_ (.A1(_2626_),
    .A2(_2736_),
    .ZN(_2794_));
 NOR2_X1 _3630_ (.A1(_2626_),
    .A2(_2736_),
    .ZN(_2795_));
 OAI21_X1 _3631_ (.A(_2794_),
    .B1(_2795_),
    .B2(_2699_),
    .ZN(_2796_));
 AND2_X1 _3632_ (.A1(_2703_),
    .A2(_2734_),
    .ZN(_2797_));
 OR2_X1 _3633_ (.A1(_2703_),
    .A2(_2734_),
    .ZN(_2798_));
 AOI21_X1 _3634_ (.A(_2797_),
    .B1(_2798_),
    .B2(_2700_),
    .ZN(_2799_));
 OR2_X1 _3635_ (.A1(_2662_),
    .A2(_2735_),
    .ZN(_2800_));
 INV_X1 _3636_ (.A(_2488_),
    .ZN(_2801_));
 NAND2_X1 _3637_ (.A1(_2519_),
    .A2(_2588_),
    .ZN(_2802_));
 OR3_X1 _3638_ (.A1(_2802_),
    .A2(_2662_),
    .A3(_2735_),
    .ZN(_2803_));
 OAI221_X1 _3639_ (.A(_2799_),
    .B1(_2800_),
    .B2(_2630_),
    .C1(_2801_),
    .C2(_2803_),
    .ZN(_2804_));
 INV_X1 _3640_ (.A(_2731_),
    .ZN(_2805_));
 NOR2_X1 _3641_ (.A1(_2805_),
    .A2(_2733_),
    .ZN(_2806_));
 NOR2_X1 _3642_ (.A1(_2704_),
    .A2(_2729_),
    .ZN(_2807_));
 AOI22_X1 _3643_ (.A1(_2657_),
    .A2(_2807_),
    .B1(_2730_),
    .B2(_0008_),
    .ZN(_2808_));
 INV_X1 _3644_ (.A(_2726_),
    .ZN(_2809_));
 NOR2_X1 _3645_ (.A1(_2716_),
    .A2(_2809_),
    .ZN(_2810_));
 NAND2_X1 _3646_ (.A1(_2718_),
    .A2(_2724_),
    .ZN(_2811_));
 NOR2_X1 _3647_ (.A1(_2718_),
    .A2(_2724_),
    .ZN(_2812_));
 OAI21_X1 _3648_ (.A(_2811_),
    .B1(_2812_),
    .B2(_2717_),
    .ZN(_2813_));
 AOI21_X1 _3649_ (.A(\iir1.y[8] ),
    .B1(\iir1.y[7] ),
    .B2(\iir1.y[9] ),
    .ZN(_2814_));
 AOI21_X1 _3650_ (.A(_2814_),
    .B1(_2574_),
    .B2(\iir1.y[7] ),
    .ZN(_2815_));
 XOR2_X1 _3651_ (.A(_2813_),
    .B(_2815_),
    .Z(_2816_));
 XOR2_X1 _3652_ (.A(_2810_),
    .B(_2816_),
    .Z(_2817_));
 AND2_X1 _3653_ (.A1(_2714_),
    .A2(_2727_),
    .ZN(_2818_));
 AOI21_X1 _3654_ (.A(_2818_),
    .B1(_2728_),
    .B2(_2712_),
    .ZN(_2819_));
 XNOR2_X1 _3655_ (.A(_2817_),
    .B(_2819_),
    .ZN(_2820_));
 XOR2_X1 _3656_ (.A(_2807_),
    .B(_2820_),
    .Z(_2821_));
 XOR2_X1 _3657_ (.A(_0030_),
    .B(_2821_),
    .Z(_2822_));
 XNOR2_X1 _3658_ (.A(_2808_),
    .B(_2822_),
    .ZN(_2823_));
 XOR2_X1 _3659_ (.A(_2806_),
    .B(_2823_),
    .Z(_2824_));
 XNOR2_X1 _3660_ (.A(_2804_),
    .B(_2824_),
    .ZN(_2825_));
 XNOR2_X1 _3661_ (.A(\iir2.x2[10] ),
    .B(_2825_),
    .ZN(_2826_));
 XOR2_X1 _3662_ (.A(_2796_),
    .B(_2826_),
    .Z(_2827_));
 XNOR2_X1 _3663_ (.A(_2793_),
    .B(_2827_),
    .ZN(_2828_));
 XNOR2_X1 _3664_ (.A(_2791_),
    .B(_2828_),
    .ZN(_2829_));
 XNOR2_X1 _3665_ (.A(_2789_),
    .B(_2829_),
    .ZN(_2830_));
 XOR2_X1 _3666_ (.A(_2788_),
    .B(_2830_),
    .Z(_2831_));
 OAI211_X1 _3667_ (.A(_2743_),
    .B(_2831_),
    .C1(_2750_),
    .C2(_2746_),
    .ZN(_2832_));
 NOR2_X1 _3668_ (.A1(_2690_),
    .A2(_2742_),
    .ZN(_2833_));
 NAND2_X1 _3669_ (.A1(_2833_),
    .A2(_2831_),
    .ZN(_2834_));
 OR2_X1 _3670_ (.A1(_2833_),
    .A2(_2831_),
    .ZN(_2835_));
 OAI211_X1 _3671_ (.A(_2832_),
    .B(_2834_),
    .C1(_2755_),
    .C2(_2835_),
    .ZN(_2836_));
 XNOR2_X1 _3672_ (.A(_2786_),
    .B(_2836_),
    .ZN(_2837_));
 XNOR2_X1 _3673_ (.A(_2760_),
    .B(_2837_),
    .ZN(_2838_));
 XNOR2_X1 _3674_ (.A(_2767_),
    .B(_2838_),
    .ZN(_2839_));
 XNOR2_X1 _3675_ (.A(_2785_),
    .B(_2839_),
    .ZN(_2840_));
 XNOR2_X1 _3676_ (.A(_2782_),
    .B(_2840_),
    .ZN(_2841_));
 XOR2_X1 _3677_ (.A(_2781_),
    .B(_2841_),
    .Z(_2842_));
 XNOR2_X1 _3678_ (.A(_2780_),
    .B(_2842_),
    .ZN(_2843_));
 NOR2_X1 _3679_ (.A1(_2779_),
    .A2(_2843_),
    .ZN(_2844_));
 XNOR2_X1 _3680_ (.A(_2779_),
    .B(_2843_),
    .ZN(_2845_));
 AND3_X1 _3681_ (.A1(_2678_),
    .A2(_2771_),
    .A3(_2772_),
    .ZN(_2846_));
 AOI21_X1 _3682_ (.A(_2678_),
    .B1(_2771_),
    .B2(_2772_),
    .ZN(_2847_));
 NOR3_X1 _3683_ (.A1(_2676_),
    .A2(_2846_),
    .A3(_2847_),
    .ZN(_2848_));
 INV_X1 _3684_ (.A(net49),
    .ZN(_2849_));
 XOR2_X1 _3685_ (.A(_2365_),
    .B(_2411_),
    .Z(_2850_));
 NAND2_X1 _3686_ (.A1(z[4]),
    .A2(_2850_),
    .ZN(_2851_));
 XNOR2_X1 _3687_ (.A(z[5]),
    .B(_2474_),
    .ZN(_2852_));
 NOR2_X1 _3688_ (.A1(_2851_),
    .A2(_2852_),
    .ZN(_2853_));
 XOR2_X1 _3689_ (.A(_2475_),
    .B(_2536_),
    .Z(_2854_));
 XNOR2_X1 _3690_ (.A(_2853_),
    .B(_2854_),
    .ZN(_2855_));
 NOR2_X1 _3691_ (.A1(_2849_),
    .A2(_2855_),
    .ZN(_2856_));
 AOI21_X1 _3692_ (.A(_2856_),
    .B1(_2854_),
    .B2(_2853_),
    .ZN(_2857_));
 XNOR2_X1 _3693_ (.A(_1330_),
    .B(_2605_),
    .ZN(_2858_));
 NOR2_X1 _3694_ (.A1(_2857_),
    .A2(_2858_),
    .ZN(_2859_));
 XOR2_X1 _3695_ (.A(_2607_),
    .B(_2675_),
    .Z(_2860_));
 AND2_X1 _3696_ (.A1(_2859_),
    .A2(_2860_),
    .ZN(_2861_));
 INV_X1 _3697_ (.A(_2861_),
    .ZN(_2862_));
 AOI21_X1 _3698_ (.A(_2677_),
    .B1(_2773_),
    .B2(_2778_),
    .ZN(_2863_));
 NOR3_X1 _3699_ (.A1(_2848_),
    .A2(_2862_),
    .A3(_2863_),
    .ZN(_2864_));
 OAI21_X1 _3700_ (.A(_2676_),
    .B1(_2846_),
    .B2(_2847_),
    .ZN(_2865_));
 AOI21_X1 _3701_ (.A(_2861_),
    .B1(_2865_),
    .B2(_2779_),
    .ZN(_2866_));
 XOR2_X1 _3702_ (.A(_2857_),
    .B(_2858_),
    .Z(_2867_));
 XOR2_X1 _3703_ (.A(_2851_),
    .B(_2852_),
    .Z(_2868_));
 XNOR2_X1 _3704_ (.A(_2406_),
    .B(_2408_),
    .ZN(_2869_));
 NAND2_X1 _3705_ (.A1(z[2]),
    .A2(_2869_),
    .ZN(_2870_));
 XOR2_X1 _3706_ (.A(_2409_),
    .B(_2410_),
    .Z(_2871_));
 XNOR2_X1 _3707_ (.A(z[3]),
    .B(_2871_),
    .ZN(_2872_));
 NOR2_X1 _3708_ (.A1(_2870_),
    .A2(_2872_),
    .ZN(_2873_));
 NAND2_X1 _3709_ (.A1(z[3]),
    .A2(_2871_),
    .ZN(_2874_));
 XNOR2_X1 _3710_ (.A(z[4]),
    .B(_2850_),
    .ZN(_2875_));
 XOR2_X1 _3711_ (.A(_2874_),
    .B(_2875_),
    .Z(_2876_));
 AND2_X1 _3712_ (.A1(_2873_),
    .A2(_2876_),
    .ZN(_2877_));
 NAND2_X1 _3713_ (.A1(_2868_),
    .A2(_2877_),
    .ZN(_2878_));
 NOR2_X1 _3714_ (.A1(_2874_),
    .A2(_2875_),
    .ZN(_2879_));
 AND2_X1 _3715_ (.A1(_2868_),
    .A2(_2879_),
    .ZN(_2880_));
 INV_X1 _3716_ (.A(_2880_),
    .ZN(_2881_));
 XNOR2_X1 _3717_ (.A(_2849_),
    .B(_2855_),
    .ZN(_2882_));
 XNOR2_X1 _3718_ (.A(_2881_),
    .B(_2882_),
    .ZN(_2883_));
 NOR2_X1 _3719_ (.A1(_2878_),
    .A2(_2883_),
    .ZN(_2884_));
 NOR2_X1 _3720_ (.A1(_2881_),
    .A2(_2882_),
    .ZN(_2885_));
 NOR2_X1 _3721_ (.A1(_2885_),
    .A2(_2884_),
    .ZN(_2886_));
 XNOR2_X1 _3722_ (.A(_2867_),
    .B(_2886_),
    .ZN(_2887_));
 XOR2_X1 _3723_ (.A(_2878_),
    .B(_2883_),
    .Z(_2888_));
 XOR2_X1 _3724_ (.A(_2404_),
    .B(_2405_),
    .Z(_2889_));
 NAND2_X1 _3725_ (.A1(z[1]),
    .A2(_2889_),
    .ZN(_2890_));
 XNOR2_X1 _3726_ (.A(z[2]),
    .B(_2869_),
    .ZN(_2891_));
 NOR2_X1 _3727_ (.A1(_2890_),
    .A2(_2891_),
    .ZN(_2892_));
 XOR2_X1 _3728_ (.A(_2870_),
    .B(_2872_),
    .Z(_2893_));
 AND2_X1 _3729_ (.A1(_2892_),
    .A2(_2893_),
    .ZN(_2894_));
 XOR2_X1 _3730_ (.A(_2873_),
    .B(_2876_),
    .Z(_2895_));
 NAND2_X1 _3731_ (.A1(_2894_),
    .A2(_2895_),
    .ZN(_2896_));
 NOR2_X1 _3732_ (.A1(_2879_),
    .A2(_2877_),
    .ZN(_2897_));
 XOR2_X1 _3733_ (.A(_2868_),
    .B(_2897_),
    .Z(_2898_));
 NOR2_X1 _3734_ (.A1(_2896_),
    .A2(_2898_),
    .ZN(_2899_));
 NAND2_X1 _3735_ (.A1(_2888_),
    .A2(_2899_),
    .ZN(_2900_));
 XNOR2_X1 _3736_ (.A(_2402_),
    .B(_2403_),
    .ZN(_2901_));
 OR2_X1 _3737_ (.A1(_2849_),
    .A2(_2901_),
    .ZN(_2902_));
 XNOR2_X1 _3738_ (.A(z[1]),
    .B(_2889_),
    .ZN(_2903_));
 NOR2_X1 _3739_ (.A1(_2902_),
    .A2(_2903_),
    .ZN(_2904_));
 XOR2_X1 _3740_ (.A(_2890_),
    .B(_2891_),
    .Z(_2905_));
 AND2_X1 _3741_ (.A1(_2904_),
    .A2(_2905_),
    .ZN(_2906_));
 XOR2_X1 _3742_ (.A(_2892_),
    .B(_2893_),
    .Z(_2907_));
 NAND2_X1 _3743_ (.A1(_2906_),
    .A2(_2907_),
    .ZN(_2908_));
 XNOR2_X1 _3744_ (.A(_2894_),
    .B(_2895_),
    .ZN(_2909_));
 OR3_X1 _3745_ (.A1(_2898_),
    .A2(_2908_),
    .A3(_2909_),
    .ZN(_2910_));
 XNOR2_X1 _3746_ (.A(_2888_),
    .B(_2899_),
    .ZN(_2911_));
 OAI21_X1 _3747_ (.A(_2900_),
    .B1(_2910_),
    .B2(_2911_),
    .ZN(_2912_));
 AOI22_X1 _3748_ (.A1(_2867_),
    .A2(_2884_),
    .B1(_2887_),
    .B2(_2912_),
    .ZN(_2913_));
 NAND2_X1 _3749_ (.A1(_2867_),
    .A2(_2885_),
    .ZN(_2914_));
 XNOR2_X1 _3750_ (.A(_2859_),
    .B(_2860_),
    .ZN(_2915_));
 XNOR2_X1 _3751_ (.A(_2914_),
    .B(_2915_),
    .ZN(_2916_));
 OR2_X1 _3752_ (.A1(_2913_),
    .A2(_2916_),
    .ZN(_2917_));
 OR3_X1 _3753_ (.A1(_2864_),
    .A2(_2866_),
    .A3(_2917_),
    .ZN(_2918_));
 OAI21_X1 _3754_ (.A(_2862_),
    .B1(_2863_),
    .B2(_2848_),
    .ZN(_2919_));
 OR2_X1 _3755_ (.A1(_2914_),
    .A2(_2915_),
    .ZN(_2920_));
 INV_X1 _3756_ (.A(_2920_),
    .ZN(_2921_));
 AOI21_X1 _3757_ (.A(_2864_),
    .B1(_2919_),
    .B2(_2921_),
    .ZN(_2922_));
 AOI21_X1 _3758_ (.A(_2845_),
    .B1(_2918_),
    .B2(_2922_),
    .ZN(_2923_));
 NOR2_X1 _3759_ (.A1(_2844_),
    .A2(_2923_),
    .ZN(_2924_));
 AND2_X1 _3760_ (.A1(_2780_),
    .A2(_2842_),
    .ZN(_2925_));
 NAND2_X1 _3761_ (.A1(_2782_),
    .A2(_2840_),
    .ZN(_2926_));
 OAI21_X1 _3762_ (.A(_2926_),
    .B1(_2841_),
    .B2(_2781_),
    .ZN(_2927_));
 NOR2_X1 _3763_ (.A1(z[4]),
    .A2(_2783_),
    .ZN(_2928_));
 INV_X1 _3764_ (.A(_2928_),
    .ZN(_2929_));
 NOR2_X1 _3765_ (.A1(_2767_),
    .A2(_2838_),
    .ZN(_2930_));
 NAND2_X1 _3766_ (.A1(_2767_),
    .A2(_2838_),
    .ZN(_2931_));
 AOI21_X1 _3767_ (.A(_2930_),
    .B1(_2931_),
    .B2(_2785_),
    .ZN(_2932_));
 NAND2_X1 _3768_ (.A1(z[4]),
    .A2(z[3]),
    .ZN(_2933_));
 NOR2_X1 _3769_ (.A1(z[5]),
    .A2(_2933_),
    .ZN(_2934_));
 OR2_X1 _3770_ (.A1(z[5]),
    .A2(z[4]),
    .ZN(_2935_));
 NAND2_X1 _3771_ (.A1(z[5]),
    .A2(z[4]),
    .ZN(_2936_));
 AOI22_X1 _3772_ (.A1(z[4]),
    .A2(z[3]),
    .B1(_2935_),
    .B2(_2936_),
    .ZN(_2937_));
 NOR2_X1 _3773_ (.A1(_2934_),
    .A2(_2937_),
    .ZN(_2938_));
 OR2_X1 _3774_ (.A1(_2760_),
    .A2(_2837_),
    .ZN(_2939_));
 NAND2_X1 _3775_ (.A1(z[10]),
    .A2(_2836_),
    .ZN(_2940_));
 NAND2_X1 _3776_ (.A1(_2743_),
    .A2(_2831_),
    .ZN(_2941_));
 AOI21_X1 _3777_ (.A(_2941_),
    .B1(_2688_),
    .B2(_2687_),
    .ZN(_2942_));
 OR2_X1 _3778_ (.A1(_2788_),
    .A2(_2830_),
    .ZN(_2943_));
 NAND2_X1 _3779_ (.A1(_2943_),
    .A2(_2834_),
    .ZN(_2944_));
 OR2_X1 _3780_ (.A1(_2791_),
    .A2(_2828_),
    .ZN(_2945_));
 OAI21_X1 _3781_ (.A(_2945_),
    .B1(_2829_),
    .B2(_2789_),
    .ZN(_2946_));
 NOR2_X1 _3782_ (.A1(_0016_),
    .A2(_2792_),
    .ZN(_2947_));
 AND2_X1 _3783_ (.A1(_2796_),
    .A2(_2826_),
    .ZN(_2948_));
 AOI21_X1 _3784_ (.A(_2948_),
    .B1(_2827_),
    .B2(_2793_),
    .ZN(_2949_));
 XOR2_X1 _3785_ (.A(\iir2.x2[10] ),
    .B(_0031_),
    .Z(_2950_));
 XNOR2_X1 _3786_ (.A(_2825_),
    .B(_2950_),
    .ZN(_2951_));
 NAND2_X1 _3787_ (.A1(_2626_),
    .A2(_2951_),
    .ZN(_0120_));
 AND2_X1 _3788_ (.A1(_2806_),
    .A2(_2823_),
    .ZN(_0121_));
 AOI21_X1 _3789_ (.A(_0121_),
    .B1(_2824_),
    .B2(_2804_),
    .ZN(_0122_));
 INV_X1 _3790_ (.A(_2808_),
    .ZN(_0123_));
 NAND2_X1 _3791_ (.A1(_0123_),
    .A2(_2822_),
    .ZN(_0124_));
 NOR2_X1 _3792_ (.A1(_2704_),
    .A2(_2820_),
    .ZN(_0125_));
 NAND2_X1 _3793_ (.A1(_2729_),
    .A2(_0125_),
    .ZN(_0126_));
 NAND2_X1 _3794_ (.A1(_0030_),
    .A2(_2821_),
    .ZN(_0127_));
 AND2_X1 _3795_ (.A1(_2813_),
    .A2(_2815_),
    .ZN(_0128_));
 OAI21_X1 _3796_ (.A(_2648_),
    .B1(_2573_),
    .B2(_2721_),
    .ZN(_0129_));
 NAND2_X1 _3797_ (.A1(\iir1.y[7] ),
    .A2(_2574_),
    .ZN(_0130_));
 OAI21_X1 _3798_ (.A(_0130_),
    .B1(_0006_),
    .B2(\iir1.y[8] ),
    .ZN(_0131_));
 XNOR2_X1 _3799_ (.A(_0129_),
    .B(_0131_),
    .ZN(_0132_));
 XNOR2_X1 _3800_ (.A(_0128_),
    .B(_0132_),
    .ZN(_0133_));
 NOR2_X1 _3801_ (.A1(_2810_),
    .A2(_2816_),
    .ZN(_0134_));
 NAND2_X1 _3802_ (.A1(_2810_),
    .A2(_2816_),
    .ZN(_0135_));
 AOI21_X1 _3803_ (.A(_0134_),
    .B1(_2819_),
    .B2(_0135_),
    .ZN(_0136_));
 XNOR2_X1 _3804_ (.A(_0133_),
    .B(_0136_),
    .ZN(_0137_));
 INV_X1 _3805_ (.A(_0004_),
    .ZN(_0138_));
 XNOR2_X1 _3806_ (.A(_0138_),
    .B(_0125_),
    .ZN(_0139_));
 XNOR2_X1 _3807_ (.A(_0137_),
    .B(_0139_),
    .ZN(_0140_));
 AND3_X1 _3808_ (.A1(_0126_),
    .A2(_0127_),
    .A3(_0140_),
    .ZN(_0141_));
 AOI21_X1 _3809_ (.A(_0140_),
    .B1(_0127_),
    .B2(_0126_),
    .ZN(_0142_));
 OR2_X1 _3810_ (.A1(_0141_),
    .A2(_0142_),
    .ZN(_0143_));
 XOR2_X1 _3811_ (.A(_0124_),
    .B(_0143_),
    .Z(_0144_));
 XNOR2_X1 _3812_ (.A(_2950_),
    .B(_0144_),
    .ZN(_0145_));
 XNOR2_X1 _3813_ (.A(_0122_),
    .B(_0145_),
    .ZN(_0146_));
 XNOR2_X1 _3814_ (.A(_0120_),
    .B(_0146_),
    .ZN(_0147_));
 XNOR2_X1 _3815_ (.A(_2698_),
    .B(_0147_),
    .ZN(_0148_));
 XOR2_X1 _3816_ (.A(_2949_),
    .B(_0148_),
    .Z(_0149_));
 XOR2_X1 _3817_ (.A(_2947_),
    .B(_0149_),
    .Z(_0150_));
 XOR2_X1 _3818_ (.A(_2946_),
    .B(_0150_),
    .Z(_0151_));
 OR3_X1 _3819_ (.A1(_2942_),
    .A2(_2944_),
    .A3(_0151_),
    .ZN(_0152_));
 OAI21_X1 _3820_ (.A(_0151_),
    .B1(_2944_),
    .B2(_2942_),
    .ZN(_0153_));
 AND2_X1 _3821_ (.A1(_0152_),
    .A2(_0153_),
    .ZN(_0154_));
 XOR2_X1 _3822_ (.A(_2940_),
    .B(_0154_),
    .Z(_0155_));
 XOR2_X1 _3823_ (.A(_2939_),
    .B(_0155_),
    .Z(_0156_));
 XNOR2_X1 _3824_ (.A(_2938_),
    .B(_0156_),
    .ZN(_0157_));
 XOR2_X1 _3825_ (.A(_2932_),
    .B(_0157_),
    .Z(_0158_));
 XNOR2_X1 _3826_ (.A(_2929_),
    .B(_0158_),
    .ZN(_0159_));
 XOR2_X1 _3827_ (.A(_2927_),
    .B(_0159_),
    .Z(_0160_));
 XOR2_X1 _3828_ (.A(_2925_),
    .B(_0160_),
    .Z(_0161_));
 XOR2_X1 _3829_ (.A(_0002_),
    .B(\iir2.y2[10] ),
    .Z(_0162_));
 XNOR2_X1 _3830_ (.A(_0161_),
    .B(_0162_),
    .ZN(_0163_));
 XNOR2_X1 _3831_ (.A(_2924_),
    .B(_0163_),
    .ZN(_0164_));
 NOR2_X1 _3832_ (.A1(_0002_),
    .A2(_0164_),
    .ZN(_0165_));
 NAND2_X1 _3833_ (.A1(_2927_),
    .A2(_0159_),
    .ZN(_0166_));
 OR2_X1 _3834_ (.A1(_2932_),
    .A2(_0157_),
    .ZN(_0167_));
 AND2_X1 _3835_ (.A1(_2932_),
    .A2(_0157_),
    .ZN(_0168_));
 OAI21_X1 _3836_ (.A(_0167_),
    .B1(_0168_),
    .B2(_2929_),
    .ZN(_0169_));
 NOR2_X1 _3837_ (.A1(_2939_),
    .A2(_0155_),
    .ZN(_0170_));
 AOI21_X1 _3838_ (.A(_0170_),
    .B1(_0156_),
    .B2(_2938_),
    .ZN(_0171_));
 XOR2_X1 _3839_ (.A(z[6]),
    .B(z[5]),
    .Z(_0172_));
 XNOR2_X1 _3840_ (.A(_2936_),
    .B(_0172_),
    .ZN(_0173_));
 INV_X1 _3841_ (.A(_0173_),
    .ZN(_0174_));
 OR2_X1 _3842_ (.A1(_2940_),
    .A2(_0154_),
    .ZN(_0175_));
 NAND2_X1 _3843_ (.A1(_2946_),
    .A2(_0150_),
    .ZN(_0176_));
 NOR2_X1 _3844_ (.A1(_2949_),
    .A2(_0148_),
    .ZN(_0177_));
 AOI21_X1 _3845_ (.A(_0177_),
    .B1(_0149_),
    .B2(_2947_),
    .ZN(_0178_));
 NOR3_X1 _3846_ (.A1(_0031_),
    .A2(_2951_),
    .A3(_0146_),
    .ZN(_0179_));
 AOI21_X1 _3847_ (.A(_0179_),
    .B1(_0147_),
    .B2(_2698_),
    .ZN(_0180_));
 AND2_X1 _3848_ (.A1(_2626_),
    .A2(_0146_),
    .ZN(_0181_));
 NAND2_X1 _3849_ (.A1(\iir1.y2[10] ),
    .A2(_0137_),
    .ZN(_0182_));
 AND2_X1 _3850_ (.A1(\iir1.y2[10] ),
    .A2(_2820_),
    .ZN(_0183_));
 OAI21_X1 _3851_ (.A(_0182_),
    .B1(_0137_),
    .B2(_0183_),
    .ZN(_0184_));
 AND2_X1 _3852_ (.A1(_0128_),
    .A2(_0132_),
    .ZN(_0185_));
 OR2_X1 _3853_ (.A1(_0128_),
    .A2(_0132_),
    .ZN(_0186_));
 AOI21_X1 _3854_ (.A(_0185_),
    .B1(_0186_),
    .B2(_0136_),
    .ZN(_0187_));
 NOR2_X1 _3855_ (.A1(_2721_),
    .A2(_2573_),
    .ZN(_0188_));
 AOI21_X1 _3856_ (.A(_0188_),
    .B1(_0131_),
    .B2(_2648_),
    .ZN(_0189_));
 NAND2_X1 _3857_ (.A1(_0187_),
    .A2(_0189_),
    .ZN(_0190_));
 NOR2_X1 _3858_ (.A1(_2704_),
    .A2(_0137_),
    .ZN(_0191_));
 XNOR2_X1 _3859_ (.A(_0004_),
    .B(_0191_),
    .ZN(_0192_));
 XNOR2_X1 _3860_ (.A(_0190_),
    .B(_0192_),
    .ZN(_0193_));
 XNOR2_X1 _3861_ (.A(_0184_),
    .B(_0193_),
    .ZN(_0194_));
 XNOR2_X1 _3862_ (.A(_0142_),
    .B(_0194_),
    .ZN(_0195_));
 NOR2_X1 _3863_ (.A1(_0124_),
    .A2(_0143_),
    .ZN(_0196_));
 AND3_X1 _3864_ (.A1(_2804_),
    .A2(_2824_),
    .A3(_0144_),
    .ZN(_0197_));
 AOI211_X1 _3865_ (.A(_0196_),
    .B(_0197_),
    .C1(_0144_),
    .C2(_0121_),
    .ZN(_0198_));
 XOR2_X1 _3866_ (.A(_0195_),
    .B(_0198_),
    .Z(_0199_));
 XNOR2_X1 _3867_ (.A(_0031_),
    .B(_0199_),
    .ZN(_0200_));
 XNOR2_X1 _3868_ (.A(_0181_),
    .B(_0200_),
    .ZN(_0201_));
 XNOR2_X1 _3869_ (.A(_0180_),
    .B(_0201_),
    .ZN(_0202_));
 XNOR2_X1 _3870_ (.A(_2792_),
    .B(_0202_),
    .ZN(_0203_));
 XOR2_X1 _3871_ (.A(_0178_),
    .B(_0203_),
    .Z(_0204_));
 INV_X1 _3872_ (.A(_0204_),
    .ZN(_0205_));
 AND3_X1 _3873_ (.A1(_0176_),
    .A2(_0153_),
    .A3(_0205_),
    .ZN(_0206_));
 AOI21_X1 _3874_ (.A(_0205_),
    .B1(_0153_),
    .B2(_0176_),
    .ZN(_0207_));
 NOR2_X1 _3875_ (.A1(_0206_),
    .A2(_0207_),
    .ZN(_0208_));
 XOR2_X1 _3876_ (.A(_0175_),
    .B(_0208_),
    .Z(_0209_));
 XNOR2_X1 _3877_ (.A(_0174_),
    .B(_0209_),
    .ZN(_0210_));
 XOR2_X1 _3878_ (.A(_0171_),
    .B(_0210_),
    .Z(_0211_));
 XOR2_X1 _3879_ (.A(_2934_),
    .B(_0211_),
    .Z(_0212_));
 XNOR2_X1 _3880_ (.A(_0169_),
    .B(_0212_),
    .ZN(_0213_));
 XOR2_X1 _3881_ (.A(_0166_),
    .B(_0213_),
    .Z(_0214_));
 INV_X1 _3882_ (.A(_0214_),
    .ZN(_0215_));
 AND2_X1 _3883_ (.A1(_2925_),
    .A2(_0160_),
    .ZN(_0216_));
 AOI21_X1 _3884_ (.A(_0216_),
    .B1(_0161_),
    .B2(_2844_),
    .ZN(_0217_));
 XNOR2_X1 _3885_ (.A(_2848_),
    .B(_2843_),
    .ZN(_0218_));
 NAND3_X1 _3886_ (.A1(_2779_),
    .A2(_2861_),
    .A3(_2865_),
    .ZN(_0219_));
 OAI21_X1 _3887_ (.A(_0219_),
    .B1(_2866_),
    .B2(_2920_),
    .ZN(_0220_));
 NOR3_X1 _3888_ (.A1(_2864_),
    .A2(_2866_),
    .A3(_2917_),
    .ZN(_0221_));
 OAI211_X1 _3889_ (.A(_0218_),
    .B(_0161_),
    .C1(_0220_),
    .C2(_0221_),
    .ZN(_0222_));
 NAND3_X1 _3890_ (.A1(_0215_),
    .A2(_0217_),
    .A3(_0222_),
    .ZN(_0223_));
 NAND2_X1 _3891_ (.A1(_2925_),
    .A2(_0160_),
    .ZN(_0224_));
 XNOR2_X1 _3892_ (.A(_2925_),
    .B(_0160_),
    .ZN(_0225_));
 OR2_X1 _3893_ (.A1(_2779_),
    .A2(_2843_),
    .ZN(_0226_));
 OAI21_X1 _3894_ (.A(_0224_),
    .B1(_0225_),
    .B2(_0226_),
    .ZN(_0227_));
 AOI211_X1 _3895_ (.A(_2845_),
    .B(_0225_),
    .C1(_2922_),
    .C2(_2918_),
    .ZN(_0228_));
 OAI21_X1 _3896_ (.A(_0214_),
    .B1(_0227_),
    .B2(_0228_),
    .ZN(_0229_));
 NAND2_X1 _3897_ (.A1(_0223_),
    .A2(_0229_),
    .ZN(_0230_));
 XNOR2_X1 _3898_ (.A(_0162_),
    .B(_0230_),
    .ZN(_0231_));
 XNOR2_X1 _3899_ (.A(_0165_),
    .B(_0231_),
    .ZN(_0232_));
 AOI21_X1 _3900_ (.A(\iir2.y2[10] ),
    .B1(_0223_),
    .B2(_0229_),
    .ZN(_0233_));
 AND3_X1 _3901_ (.A1(\iir2.y2[10] ),
    .A2(_0223_),
    .A3(_0229_),
    .ZN(_0234_));
 NOR3_X1 _3902_ (.A1(_0002_),
    .A2(_0233_),
    .A3(_0234_),
    .ZN(_0235_));
 AOI22_X1 _3903_ (.A1(_1319_),
    .A2(_0232_),
    .B1(_0235_),
    .B2(_0164_),
    .ZN(_0236_));
 XOR2_X1 _3904_ (.A(\iir2.y2[10] ),
    .B(\iir2.y2[9] ),
    .Z(_0237_));
 NOR2_X1 _3905_ (.A1(_0166_),
    .A2(_0213_),
    .ZN(_0238_));
 AOI21_X1 _3906_ (.A(_0215_),
    .B1(_0217_),
    .B2(_0222_),
    .ZN(_0239_));
 NOR2_X1 _3907_ (.A1(_0238_),
    .A2(_0239_),
    .ZN(_0240_));
 NAND2_X1 _3908_ (.A1(_0169_),
    .A2(_0212_),
    .ZN(_0241_));
 NOR2_X1 _3909_ (.A1(_0171_),
    .A2(_0210_),
    .ZN(_0242_));
 AOI21_X1 _3910_ (.A(_0242_),
    .B1(_0211_),
    .B2(_2934_),
    .ZN(_0243_));
 NOR2_X1 _3911_ (.A1(z[6]),
    .A2(_2936_),
    .ZN(_0244_));
 AOI21_X1 _3912_ (.A(_2786_),
    .B1(_0152_),
    .B2(_0153_),
    .ZN(_0245_));
 OAI21_X1 _3913_ (.A(_0245_),
    .B1(_0207_),
    .B2(_0206_),
    .ZN(_0246_));
 OAI22_X1 _3914_ (.A1(_0174_),
    .A2(_0209_),
    .B1(_0246_),
    .B2(_2836_),
    .ZN(_0247_));
 NAND2_X1 _3915_ (.A1(z[6]),
    .A2(z[5]),
    .ZN(_0248_));
 NOR2_X1 _3916_ (.A1(z[7]),
    .A2(_0248_),
    .ZN(_0249_));
 OR2_X1 _3917_ (.A1(z[7]),
    .A2(z[6]),
    .ZN(_0250_));
 NAND2_X1 _3918_ (.A1(z[7]),
    .A2(z[6]),
    .ZN(_0251_));
 AOI22_X1 _3919_ (.A1(z[6]),
    .A2(z[5]),
    .B1(_0250_),
    .B2(_0251_),
    .ZN(_0252_));
 NOR2_X1 _3920_ (.A1(_0249_),
    .A2(_0252_),
    .ZN(_0253_));
 OR2_X1 _3921_ (.A1(_0178_),
    .A2(_0203_),
    .ZN(_0254_));
 OAI21_X1 _3922_ (.A(_0254_),
    .B1(_0205_),
    .B2(_0176_),
    .ZN(_0255_));
 NAND2_X1 _3923_ (.A1(_0151_),
    .A2(_0204_),
    .ZN(_0256_));
 AOI21_X1 _3924_ (.A(_0256_),
    .B1(_2834_),
    .B2(_2943_),
    .ZN(_0257_));
 NAND4_X1 _3925_ (.A1(_2743_),
    .A2(_2831_),
    .A3(_0151_),
    .A4(_0204_),
    .ZN(_0258_));
 NAND3_X1 _3926_ (.A1(_2541_),
    .A2(_2601_),
    .A3(_2670_),
    .ZN(_0259_));
 AOI21_X1 _3927_ (.A(_0258_),
    .B1(_0259_),
    .B2(_2687_),
    .ZN(_0260_));
 NOR2_X1 _3928_ (.A1(_2473_),
    .A2(_2532_),
    .ZN(_0261_));
 NAND3_X1 _3929_ (.A1(_0261_),
    .A2(_2601_),
    .A3(_2670_),
    .ZN(_0262_));
 NOR3_X1 _3930_ (.A1(_2412_),
    .A2(_0262_),
    .A3(_0258_),
    .ZN(_0263_));
 NOR4_X1 _3931_ (.A1(_0255_),
    .A2(_0257_),
    .A3(_0260_),
    .A4(_0263_),
    .ZN(_0264_));
 OR2_X1 _3932_ (.A1(_0180_),
    .A2(_0201_),
    .ZN(_0265_));
 OAI21_X1 _3933_ (.A(_0265_),
    .B1(_0202_),
    .B2(_2792_),
    .ZN(_0266_));
 AND2_X1 _3934_ (.A1(_0181_),
    .A2(_0200_),
    .ZN(_0267_));
 AND2_X1 _3935_ (.A1(_2626_),
    .A2(_0199_),
    .ZN(_0268_));
 NAND2_X1 _3936_ (.A1(_0142_),
    .A2(_0194_),
    .ZN(_0269_));
 OAI21_X1 _3937_ (.A(_0269_),
    .B1(_0195_),
    .B2(_0198_),
    .ZN(_0270_));
 OAI211_X1 _3938_ (.A(_0182_),
    .B(_0193_),
    .C1(_0183_),
    .C2(_0137_),
    .ZN(_0271_));
 MUX2_X1 _3939_ (.A(_0182_),
    .B(\iir1.y2[10] ),
    .S(_0190_),
    .Z(_0272_));
 INV_X1 _3940_ (.A(_0272_),
    .ZN(_0273_));
 NOR2_X1 _3941_ (.A1(_2704_),
    .A2(_0190_),
    .ZN(_0274_));
 XNOR2_X1 _3942_ (.A(\iir1.y[10] ),
    .B(_0004_),
    .ZN(_0275_));
 XNOR2_X1 _3943_ (.A(_0274_),
    .B(_0275_),
    .ZN(_0276_));
 XNOR2_X1 _3944_ (.A(_0273_),
    .B(_0276_),
    .ZN(_0277_));
 XOR2_X1 _3945_ (.A(_0271_),
    .B(_0277_),
    .Z(_0278_));
 XNOR2_X1 _3946_ (.A(_0270_),
    .B(_0278_),
    .ZN(_0279_));
 XNOR2_X1 _3947_ (.A(_2626_),
    .B(_0279_),
    .ZN(_0280_));
 XOR2_X1 _3948_ (.A(_0268_),
    .B(_0280_),
    .Z(_0281_));
 XNOR2_X1 _3949_ (.A(_0267_),
    .B(_0281_),
    .ZN(_0282_));
 XNOR2_X1 _3950_ (.A(\iir2.x2[10] ),
    .B(_0282_),
    .ZN(_0283_));
 XNOR2_X1 _3951_ (.A(_0266_),
    .B(_0283_),
    .ZN(_0284_));
 XOR2_X1 _3952_ (.A(_0264_),
    .B(_0284_),
    .Z(_0285_));
 XNOR2_X1 _3953_ (.A(_0246_),
    .B(_0285_),
    .ZN(_0286_));
 XOR2_X1 _3954_ (.A(_0253_),
    .B(_0286_),
    .Z(_0287_));
 XNOR2_X1 _3955_ (.A(_0247_),
    .B(_0287_),
    .ZN(_0288_));
 XNOR2_X1 _3956_ (.A(_0244_),
    .B(_0288_),
    .ZN(_0289_));
 XOR2_X1 _3957_ (.A(_0243_),
    .B(_0289_),
    .Z(_0290_));
 XOR2_X1 _3958_ (.A(_0241_),
    .B(_0290_),
    .Z(_0291_));
 XNOR2_X1 _3959_ (.A(_0162_),
    .B(_0291_),
    .ZN(_0292_));
 XNOR2_X1 _3960_ (.A(_0240_),
    .B(_0292_),
    .ZN(_0293_));
 XOR2_X1 _3961_ (.A(_0235_),
    .B(_0293_),
    .Z(_0294_));
 XNOR2_X1 _3962_ (.A(_0237_),
    .B(_0294_),
    .ZN(_0295_));
 NOR2_X1 _3963_ (.A1(_0236_),
    .A2(_0295_),
    .ZN(_0296_));
 INV_X1 _3964_ (.A(\iir2.y2[6] ),
    .ZN(_0297_));
 NAND2_X1 _3965_ (.A1(\iir2.y2[10] ),
    .A2(\iir2.y2[8] ),
    .ZN(_0298_));
 XNOR2_X1 _3966_ (.A(_0297_),
    .B(_0298_),
    .ZN(_0299_));
 XOR2_X1 _3967_ (.A(_0236_),
    .B(_0295_),
    .Z(_0300_));
 AOI21_X1 _3968_ (.A(_0296_),
    .B1(_0299_),
    .B2(_0300_),
    .ZN(_0301_));
 NAND2_X1 _3969_ (.A1(\iir2.y2[10] ),
    .A2(\iir2.y2[9] ),
    .ZN(_0302_));
 XOR2_X1 _3970_ (.A(\iir2.y2[7] ),
    .B(_0302_),
    .Z(_0303_));
 NOR3_X1 _3971_ (.A1(_0002_),
    .A2(_0231_),
    .A3(_0293_),
    .ZN(_0304_));
 AOI21_X1 _3972_ (.A(_0304_),
    .B1(_0294_),
    .B2(_0237_),
    .ZN(_0305_));
 NOR2_X1 _3973_ (.A1(_0002_),
    .A2(_0293_),
    .ZN(_0306_));
 INV_X1 _3974_ (.A(_0243_),
    .ZN(_0307_));
 NAND2_X1 _3975_ (.A1(_0307_),
    .A2(_0289_),
    .ZN(_0308_));
 AND2_X1 _3976_ (.A1(_0247_),
    .A2(_0287_),
    .ZN(_0309_));
 NOR3_X1 _3977_ (.A1(z[6]),
    .A2(_2936_),
    .A3(_0288_),
    .ZN(_0310_));
 NOR3_X1 _3978_ (.A1(_2786_),
    .A2(_0208_),
    .A3(_0285_),
    .ZN(_0311_));
 AOI22_X1 _3979_ (.A1(_0253_),
    .A2(_0286_),
    .B1(_0311_),
    .B2(_0154_),
    .ZN(_0312_));
 NOR2_X1 _3980_ (.A1(z[8]),
    .A2(_0251_),
    .ZN(_0313_));
 OR2_X1 _3981_ (.A1(z[8]),
    .A2(z[7]),
    .ZN(_0314_));
 NAND2_X1 _3982_ (.A1(z[8]),
    .A2(z[7]),
    .ZN(_0315_));
 AOI22_X1 _3983_ (.A1(z[7]),
    .A2(z[6]),
    .B1(_0314_),
    .B2(_0315_),
    .ZN(_0316_));
 NOR2_X1 _3984_ (.A1(_0313_),
    .A2(_0316_),
    .ZN(_0317_));
 XNOR2_X1 _3985_ (.A(_0264_),
    .B(_0284_),
    .ZN(_0318_));
 OAI211_X1 _3986_ (.A(z[10]),
    .B(_0318_),
    .C1(_0207_),
    .C2(_0206_),
    .ZN(_0319_));
 NAND2_X1 _3987_ (.A1(_0266_),
    .A2(_0283_),
    .ZN(_0320_));
 OAI21_X1 _3988_ (.A(_0320_),
    .B1(_0284_),
    .B2(_0264_),
    .ZN(_0321_));
 NOR2_X1 _3989_ (.A1(_2554_),
    .A2(_0282_),
    .ZN(_0322_));
 AOI21_X1 _3990_ (.A(_0322_),
    .B1(_0281_),
    .B2(_0267_),
    .ZN(_0323_));
 NAND2_X1 _3991_ (.A1(_0279_),
    .A2(_0268_),
    .ZN(_0324_));
 NOR2_X1 _3992_ (.A1(_0031_),
    .A2(_0279_),
    .ZN(_0325_));
 NOR2_X1 _3993_ (.A1(_0271_),
    .A2(_0277_),
    .ZN(_0326_));
 AOI21_X1 _3994_ (.A(_0326_),
    .B1(_0278_),
    .B2(_0270_),
    .ZN(_0327_));
 NAND2_X1 _3995_ (.A1(_0273_),
    .A2(_0276_),
    .ZN(_0328_));
 AOI21_X1 _3996_ (.A(_2704_),
    .B1(_0187_),
    .B2(_0189_),
    .ZN(_0329_));
 MUX2_X1 _3997_ (.A(_0329_),
    .B(_2704_),
    .S(\iir1.y[10] ),
    .Z(_0330_));
 NOR2_X1 _3998_ (.A1(\iir1.y2[10] ),
    .A2(\iir1.y[10] ),
    .ZN(_0331_));
 XNOR2_X1 _3999_ (.A(_0004_),
    .B(_0331_),
    .ZN(_0332_));
 XOR2_X1 _4000_ (.A(_0330_),
    .B(_0332_),
    .Z(_0333_));
 XNOR2_X1 _4001_ (.A(_0328_),
    .B(_0333_),
    .ZN(_0334_));
 XOR2_X1 _4002_ (.A(_0327_),
    .B(_0334_),
    .Z(_0335_));
 XNOR2_X1 _4003_ (.A(_2626_),
    .B(_0335_),
    .ZN(_0336_));
 XNOR2_X1 _4004_ (.A(_0325_),
    .B(_0336_),
    .ZN(_0337_));
 XOR2_X1 _4005_ (.A(_0324_),
    .B(_0337_),
    .Z(_0338_));
 XNOR2_X1 _4006_ (.A(\iir2.x2[10] ),
    .B(_0338_),
    .ZN(_0339_));
 XOR2_X1 _4007_ (.A(_0323_),
    .B(_0339_),
    .Z(_0340_));
 XNOR2_X1 _4008_ (.A(_0321_),
    .B(_0340_),
    .ZN(_0341_));
 XOR2_X1 _4009_ (.A(_0319_),
    .B(_0341_),
    .Z(_0342_));
 XNOR2_X1 _4010_ (.A(_0317_),
    .B(_0342_),
    .ZN(_0343_));
 XOR2_X1 _4011_ (.A(_0312_),
    .B(_0343_),
    .Z(_0344_));
 XOR2_X1 _4012_ (.A(_0249_),
    .B(_0344_),
    .Z(_0345_));
 OR3_X1 _4013_ (.A1(_0309_),
    .A2(_0310_),
    .A3(_0345_),
    .ZN(_0346_));
 OAI21_X1 _4014_ (.A(_0345_),
    .B1(_0310_),
    .B2(_0309_),
    .ZN(_0347_));
 NAND2_X1 _4015_ (.A1(_0346_),
    .A2(_0347_),
    .ZN(_0348_));
 XOR2_X1 _4016_ (.A(_0308_),
    .B(_0348_),
    .Z(_0349_));
 NAND2_X1 _4017_ (.A1(_0214_),
    .A2(_0291_),
    .ZN(_0350_));
 AOI21_X1 _4018_ (.A(_0350_),
    .B1(_0222_),
    .B2(_0217_),
    .ZN(_0351_));
 NAND2_X1 _4019_ (.A1(_0238_),
    .A2(_0291_),
    .ZN(_0352_));
 OAI21_X1 _4020_ (.A(_0352_),
    .B1(_0290_),
    .B2(_0241_),
    .ZN(_0353_));
 OR3_X1 _4021_ (.A1(_0349_),
    .A2(_0351_),
    .A3(_0353_),
    .ZN(_0354_));
 OAI21_X1 _4022_ (.A(_0349_),
    .B1(_0351_),
    .B2(_0353_),
    .ZN(_0355_));
 AND2_X1 _4023_ (.A1(_0354_),
    .A2(_0355_),
    .ZN(_0356_));
 XNOR2_X1 _4024_ (.A(_0162_),
    .B(_0356_),
    .ZN(_0357_));
 XNOR2_X1 _4025_ (.A(_0306_),
    .B(_0357_),
    .ZN(_0358_));
 XOR2_X1 _4026_ (.A(_0305_),
    .B(_0358_),
    .Z(_0359_));
 XNOR2_X1 _4027_ (.A(_0303_),
    .B(_0359_),
    .ZN(_0360_));
 NOR2_X1 _4028_ (.A1(_0301_),
    .A2(_0360_),
    .ZN(_0361_));
 XOR2_X1 _4029_ (.A(_0301_),
    .B(_0360_),
    .Z(_0362_));
 NOR2_X1 _4030_ (.A1(\iir2.y2[6] ),
    .A2(_0298_),
    .ZN(_0363_));
 AOI21_X1 _4031_ (.A(_0361_),
    .B1(_0362_),
    .B2(_0363_),
    .ZN(_0364_));
 INV_X1 _4032_ (.A(_0364_),
    .ZN(_0365_));
 NOR2_X1 _4033_ (.A1(\iir2.y2[7] ),
    .A2(_0302_),
    .ZN(_0366_));
 NOR2_X1 _4034_ (.A1(_0305_),
    .A2(_0358_),
    .ZN(_0367_));
 AOI21_X1 _4035_ (.A(_0367_),
    .B1(_0359_),
    .B2(_0303_),
    .ZN(_0368_));
 NOR3_X1 _4036_ (.A1(_0002_),
    .A2(_0293_),
    .A3(_0357_),
    .ZN(_0369_));
 NOR2_X1 _4037_ (.A1(_0308_),
    .A2(_0348_),
    .ZN(_0370_));
 INV_X1 _4038_ (.A(_0370_),
    .ZN(_0371_));
 OR2_X1 _4039_ (.A1(_0312_),
    .A2(_0343_),
    .ZN(_0372_));
 NAND2_X1 _4040_ (.A1(_0249_),
    .A2(_0344_),
    .ZN(_0373_));
 NAND2_X1 _4041_ (.A1(_0372_),
    .A2(_0373_),
    .ZN(_0374_));
 NAND3_X1 _4042_ (.A1(z[10]),
    .A2(_0318_),
    .A3(_0341_),
    .ZN(_0375_));
 INV_X1 _4043_ (.A(_0375_),
    .ZN(_0376_));
 AOI22_X1 _4044_ (.A1(_0317_),
    .A2(_0342_),
    .B1(_0376_),
    .B2(_0208_),
    .ZN(_0377_));
 XOR2_X1 _4045_ (.A(z[9]),
    .B(z[8]),
    .Z(_0378_));
 XNOR2_X1 _4046_ (.A(_0315_),
    .B(_0378_),
    .ZN(_0379_));
 NOR2_X1 _4047_ (.A1(_0323_),
    .A2(_0339_),
    .ZN(_0380_));
 AOI21_X1 _4048_ (.A(_0380_),
    .B1(_0340_),
    .B2(_0321_),
    .ZN(_0381_));
 NAND2_X1 _4049_ (.A1(\iir2.x2[10] ),
    .A2(_0338_),
    .ZN(_0382_));
 OAI21_X1 _4050_ (.A(_0382_),
    .B1(_0337_),
    .B2(_0324_),
    .ZN(_0383_));
 AND2_X1 _4051_ (.A1(_0325_),
    .A2(_0335_),
    .ZN(_0384_));
 NOR2_X1 _4052_ (.A1(_0031_),
    .A2(_0335_),
    .ZN(_0385_));
 INV_X1 _4053_ (.A(_0327_),
    .ZN(_0386_));
 NAND2_X1 _4054_ (.A1(_0386_),
    .A2(_0334_),
    .ZN(_0387_));
 AND3_X1 _4055_ (.A1(\iir1.y2[10] ),
    .A2(\iir1.y[10] ),
    .A3(_0004_),
    .ZN(_0388_));
 AOI21_X1 _4056_ (.A(_0388_),
    .B1(_0332_),
    .B2(_0330_),
    .ZN(_0389_));
 INV_X1 _4057_ (.A(_0333_),
    .ZN(_0390_));
 OAI211_X1 _4058_ (.A(_0387_),
    .B(_0389_),
    .C1(_0328_),
    .C2(_0390_),
    .ZN(_0391_));
 XNOR2_X1 _4059_ (.A(\iir2.x2[10] ),
    .B(_0391_),
    .ZN(_0392_));
 XOR2_X1 _4060_ (.A(_0385_),
    .B(_0392_),
    .Z(_0393_));
 NOR2_X1 _4061_ (.A1(_0384_),
    .A2(_0393_),
    .ZN(_0394_));
 NAND2_X1 _4062_ (.A1(_0384_),
    .A2(_0392_),
    .ZN(_0395_));
 INV_X1 _4063_ (.A(_0395_),
    .ZN(_0396_));
 NOR2_X1 _4064_ (.A1(_0394_),
    .A2(_0396_),
    .ZN(_0397_));
 XNOR2_X1 _4065_ (.A(_2554_),
    .B(_0397_),
    .ZN(_0398_));
 XOR2_X1 _4066_ (.A(_0383_),
    .B(_0398_),
    .Z(_0399_));
 XOR2_X1 _4067_ (.A(_0381_),
    .B(_0399_),
    .Z(_0400_));
 XOR2_X1 _4068_ (.A(_0375_),
    .B(_0400_),
    .Z(_0401_));
 XOR2_X1 _4069_ (.A(_0379_),
    .B(_0401_),
    .Z(_0402_));
 XOR2_X1 _4070_ (.A(_0377_),
    .B(_0402_),
    .Z(_0403_));
 XOR2_X1 _4071_ (.A(_0313_),
    .B(_0403_),
    .Z(_0404_));
 XOR2_X1 _4072_ (.A(_0374_),
    .B(_0404_),
    .Z(_0405_));
 XOR2_X1 _4073_ (.A(_0347_),
    .B(_0405_),
    .Z(_0406_));
 INV_X1 _4074_ (.A(_0406_),
    .ZN(_0407_));
 AND3_X1 _4075_ (.A1(_0371_),
    .A2(_0355_),
    .A3(_0407_),
    .ZN(_0408_));
 AOI21_X1 _4076_ (.A(_0407_),
    .B1(_0355_),
    .B2(_0371_),
    .ZN(_0409_));
 NOR2_X1 _4077_ (.A1(_0408_),
    .A2(_0409_),
    .ZN(_0410_));
 XNOR2_X1 _4078_ (.A(_0162_),
    .B(_0410_),
    .ZN(_0411_));
 XOR2_X1 _4079_ (.A(_0369_),
    .B(_0411_),
    .Z(_0412_));
 XNOR2_X1 _4080_ (.A(_1308_),
    .B(_0412_),
    .ZN(_0413_));
 XOR2_X1 _4081_ (.A(_0368_),
    .B(_0413_),
    .Z(_0414_));
 XOR2_X1 _4082_ (.A(_0366_),
    .B(_0414_),
    .Z(_0415_));
 AND2_X1 _4083_ (.A1(_0365_),
    .A2(_0415_),
    .ZN(_0416_));
 NOR3_X1 _4084_ (.A1(_0220_),
    .A2(_0221_),
    .A3(_0218_),
    .ZN(_0417_));
 NOR2_X1 _4085_ (.A1(_2923_),
    .A2(_0417_),
    .ZN(_0418_));
 XNOR2_X1 _4086_ (.A(_0162_),
    .B(_0418_),
    .ZN(_0419_));
 NOR2_X1 _4087_ (.A1(_0002_),
    .A2(_0419_),
    .ZN(_0420_));
 XOR2_X1 _4088_ (.A(_0164_),
    .B(_0420_),
    .Z(_0421_));
 XOR2_X1 _4089_ (.A(\iir2.y2[10] ),
    .B(\iir2.y2[7] ),
    .Z(_0422_));
 AOI22_X1 _4090_ (.A1(_0165_),
    .A2(_0419_),
    .B1(_0421_),
    .B2(_0422_),
    .ZN(_0423_));
 XNOR2_X1 _4091_ (.A(_1319_),
    .B(_0232_),
    .ZN(_0424_));
 NOR2_X1 _4092_ (.A1(_0423_),
    .A2(_0424_),
    .ZN(_0425_));
 INV_X1 _4093_ (.A(\iir2.y2[5] ),
    .ZN(_0426_));
 NAND2_X1 _4094_ (.A1(\iir2.y2[10] ),
    .A2(\iir2.y2[7] ),
    .ZN(_0427_));
 XNOR2_X1 _4095_ (.A(_0426_),
    .B(_0427_),
    .ZN(_0428_));
 XOR2_X1 _4096_ (.A(_0423_),
    .B(_0424_),
    .Z(_0429_));
 AOI21_X1 _4097_ (.A(_0425_),
    .B1(_0428_),
    .B2(_0429_),
    .ZN(_0430_));
 XNOR2_X1 _4098_ (.A(_0299_),
    .B(_0300_),
    .ZN(_0431_));
 NOR2_X1 _4099_ (.A1(_0430_),
    .A2(_0431_),
    .ZN(_0432_));
 XOR2_X1 _4100_ (.A(_0430_),
    .B(_0431_),
    .Z(_0433_));
 NOR2_X1 _4101_ (.A1(\iir2.y2[5] ),
    .A2(_0427_),
    .ZN(_0434_));
 AOI21_X1 _4102_ (.A(_0432_),
    .B1(_0433_),
    .B2(_0434_),
    .ZN(_0435_));
 XOR2_X1 _4103_ (.A(_0363_),
    .B(_0362_),
    .Z(_0436_));
 INV_X1 _4104_ (.A(_0436_),
    .ZN(_0437_));
 NOR2_X1 _4105_ (.A1(_0435_),
    .A2(_0437_),
    .ZN(_0438_));
 XNOR2_X1 _4106_ (.A(_0435_),
    .B(_0436_),
    .ZN(_0439_));
 INV_X1 _4107_ (.A(\iir2.y2[10] ),
    .ZN(_0440_));
 OAI21_X1 _4108_ (.A(_0440_),
    .B1(_2923_),
    .B2(_0417_),
    .ZN(_0441_));
 OR3_X1 _4109_ (.A1(_0440_),
    .A2(_2923_),
    .A3(_0417_),
    .ZN(_0442_));
 OAI21_X1 _4110_ (.A(_2920_),
    .B1(_2913_),
    .B2(_2916_),
    .ZN(_0443_));
 AOI21_X1 _4111_ (.A(_0443_),
    .B1(_2919_),
    .B2(_0219_),
    .ZN(_0444_));
 AND3_X1 _4112_ (.A1(_0219_),
    .A2(_2919_),
    .A3(_0443_),
    .ZN(_0445_));
 NOR3_X1 _4113_ (.A1(_0002_),
    .A2(_0444_),
    .A3(_0445_),
    .ZN(_0446_));
 XNOR2_X1 _4114_ (.A(\iir2.y2[10] ),
    .B(\iir2.y2[9] ),
    .ZN(_0447_));
 INV_X1 _4115_ (.A(_0002_),
    .ZN(_0448_));
 OAI211_X1 _4116_ (.A(_2920_),
    .B(_2917_),
    .C1(_2864_),
    .C2(_2866_),
    .ZN(_0449_));
 NAND3_X1 _4117_ (.A1(_0219_),
    .A2(_2919_),
    .A3(_0443_),
    .ZN(_0450_));
 AOI21_X1 _4118_ (.A(_0448_),
    .B1(_0449_),
    .B2(_0450_),
    .ZN(_0451_));
 NOR3_X1 _4119_ (.A1(_0447_),
    .A2(_0446_),
    .A3(_0451_),
    .ZN(_0452_));
 OAI211_X1 _4120_ (.A(_0441_),
    .B(_0442_),
    .C1(_0446_),
    .C2(_0452_),
    .ZN(_0453_));
 XOR2_X1 _4121_ (.A(_0026_),
    .B(_0302_),
    .Z(_0454_));
 NAND3_X1 _4122_ (.A1(_0448_),
    .A2(_0449_),
    .A3(_0450_),
    .ZN(_0455_));
 OAI21_X1 _4123_ (.A(_0002_),
    .B1(_0444_),
    .B2(_0445_),
    .ZN(_0456_));
 NAND3_X1 _4124_ (.A1(_0237_),
    .A2(_0455_),
    .A3(_0456_),
    .ZN(_0457_));
 AND4_X1 _4125_ (.A1(_0441_),
    .A2(_0442_),
    .A3(_0455_),
    .A4(_0457_),
    .ZN(_0458_));
 AOI22_X1 _4126_ (.A1(_0441_),
    .A2(_0442_),
    .B1(_0455_),
    .B2(_0457_),
    .ZN(_0459_));
 OAI21_X1 _4127_ (.A(_0454_),
    .B1(_0458_),
    .B2(_0459_),
    .ZN(_0460_));
 AND2_X1 _4128_ (.A1(_0453_),
    .A2(_0460_),
    .ZN(_0461_));
 XNOR2_X1 _4129_ (.A(_0422_),
    .B(_0421_),
    .ZN(_0462_));
 NOR2_X1 _4130_ (.A1(_0461_),
    .A2(_0462_),
    .ZN(_0463_));
 NOR2_X1 _4131_ (.A1(_0026_),
    .A2(_0302_),
    .ZN(_0464_));
 XNOR2_X1 _4132_ (.A(\iir2.y2[4] ),
    .B(_0464_),
    .ZN(_0465_));
 XOR2_X1 _4133_ (.A(_0461_),
    .B(_0462_),
    .Z(_0466_));
 AOI21_X1 _4134_ (.A(_0463_),
    .B1(_0465_),
    .B2(_0466_),
    .ZN(_0467_));
 XNOR2_X1 _4135_ (.A(_0428_),
    .B(_0429_),
    .ZN(_0468_));
 NOR2_X1 _4136_ (.A1(_0467_),
    .A2(_0468_),
    .ZN(_0469_));
 XOR2_X1 _4137_ (.A(_0467_),
    .B(_0468_),
    .Z(_0470_));
 NOR3_X1 _4138_ (.A1(\iir2.y2[4] ),
    .A2(_0026_),
    .A3(_0302_),
    .ZN(_0471_));
 AOI21_X1 _4139_ (.A(_0469_),
    .B1(_0470_),
    .B2(_0471_),
    .ZN(_0472_));
 XNOR2_X1 _4140_ (.A(_0434_),
    .B(_0433_),
    .ZN(_0473_));
 NOR2_X1 _4141_ (.A1(_0472_),
    .A2(_0473_),
    .ZN(_0474_));
 AOI21_X1 _4142_ (.A(_0438_),
    .B1(_0439_),
    .B2(_0474_),
    .ZN(_0475_));
 XOR2_X1 _4143_ (.A(_0472_),
    .B(_0473_),
    .Z(_0476_));
 NAND2_X1 _4144_ (.A1(_0439_),
    .A2(_0476_),
    .ZN(_0477_));
 XOR2_X1 _4145_ (.A(_2887_),
    .B(_2912_),
    .Z(_0478_));
 OR2_X1 _4146_ (.A1(\iir2.y2[10] ),
    .A2(_0478_),
    .ZN(_0479_));
 XOR2_X1 _4147_ (.A(_2913_),
    .B(_2916_),
    .Z(_0480_));
 XNOR2_X1 _4148_ (.A(_0162_),
    .B(_0480_),
    .ZN(_0481_));
 NAND2_X1 _4149_ (.A1(_0479_),
    .A2(_0481_),
    .ZN(_0482_));
 XOR2_X1 _4150_ (.A(\iir2.y2[9] ),
    .B(\iir2.y2[8] ),
    .Z(_0483_));
 INV_X1 _4151_ (.A(_0483_),
    .ZN(_0484_));
 NOR2_X1 _4152_ (.A1(_0479_),
    .A2(_0481_),
    .ZN(_0485_));
 OAI21_X1 _4153_ (.A(_0482_),
    .B1(_0484_),
    .B2(_0485_),
    .ZN(_0486_));
 OAI21_X1 _4154_ (.A(_0447_),
    .B1(_0446_),
    .B2(_0451_),
    .ZN(_0487_));
 NAND3_X1 _4155_ (.A1(_0457_),
    .A2(_0486_),
    .A3(_0487_),
    .ZN(_0488_));
 NAND2_X1 _4156_ (.A1(\iir2.y2[9] ),
    .A2(\iir2.y2[8] ),
    .ZN(_0489_));
 XNOR2_X1 _4157_ (.A(_0028_),
    .B(_0489_),
    .ZN(_0490_));
 AOI21_X1 _4158_ (.A(_0486_),
    .B1(_0487_),
    .B2(_0457_),
    .ZN(_0491_));
 OAI21_X1 _4159_ (.A(_0488_),
    .B1(_0490_),
    .B2(_0491_),
    .ZN(_0492_));
 OR3_X1 _4160_ (.A1(_0454_),
    .A2(_0458_),
    .A3(_0459_),
    .ZN(_0493_));
 AND3_X1 _4161_ (.A1(_0460_),
    .A2(_0492_),
    .A3(_0493_),
    .ZN(_0494_));
 INV_X1 _4162_ (.A(_0494_),
    .ZN(_0495_));
 INV_X1 _4163_ (.A(\iir2.y2[3] ),
    .ZN(_0496_));
 NOR2_X1 _4164_ (.A1(_0028_),
    .A2(_0489_),
    .ZN(_0497_));
 XNOR2_X1 _4165_ (.A(_0496_),
    .B(_0497_),
    .ZN(_0498_));
 AOI21_X1 _4166_ (.A(_0492_),
    .B1(_0493_),
    .B2(_0460_),
    .ZN(_0499_));
 OR3_X1 _4167_ (.A1(_0494_),
    .A2(_0498_),
    .A3(_0499_),
    .ZN(_0500_));
 AND2_X1 _4168_ (.A1(_0495_),
    .A2(_0500_),
    .ZN(_0501_));
 XNOR2_X1 _4169_ (.A(_0465_),
    .B(_0466_),
    .ZN(_0502_));
 NOR2_X1 _4170_ (.A1(_0501_),
    .A2(_0502_),
    .ZN(_0503_));
 XOR2_X1 _4171_ (.A(_0501_),
    .B(_0502_),
    .Z(_0504_));
 NOR3_X1 _4172_ (.A1(\iir2.y2[3] ),
    .A2(_0028_),
    .A3(_0489_),
    .ZN(_0505_));
 AOI21_X1 _4173_ (.A(_0503_),
    .B1(_0504_),
    .B2(_0505_),
    .ZN(_0506_));
 XNOR2_X1 _4174_ (.A(_0471_),
    .B(_0470_),
    .ZN(_0507_));
 NOR2_X1 _4175_ (.A1(_0506_),
    .A2(_0507_),
    .ZN(_0508_));
 XOR2_X1 _4176_ (.A(_0506_),
    .B(_0507_),
    .Z(_0509_));
 XOR2_X1 _4177_ (.A(_0479_),
    .B(_0481_),
    .Z(_0510_));
 AOI22_X1 _4178_ (.A1(_0479_),
    .A2(_0481_),
    .B1(_0483_),
    .B2(_0510_),
    .ZN(_0511_));
 AOI21_X1 _4179_ (.A(_0237_),
    .B1(_0455_),
    .B2(_0456_),
    .ZN(_0512_));
 NOR3_X1 _4180_ (.A1(_0452_),
    .A2(_0511_),
    .A3(_0512_),
    .ZN(_0513_));
 NOR3_X1 _4181_ (.A1(_0513_),
    .A2(_0490_),
    .A3(_0491_),
    .ZN(_0514_));
 XOR2_X1 _4182_ (.A(_2910_),
    .B(_2911_),
    .Z(_0515_));
 NAND2_X1 _4183_ (.A1(\iir2.y2[9] ),
    .A2(_0515_),
    .ZN(_0516_));
 XNOR2_X1 _4184_ (.A(\iir2.y2[9] ),
    .B(_0515_),
    .ZN(_0517_));
 INV_X1 _4185_ (.A(\iir2.y2[8] ),
    .ZN(_0518_));
 OAI21_X1 _4186_ (.A(_0516_),
    .B1(_0517_),
    .B2(_0518_),
    .ZN(_0519_));
 INV_X1 _4187_ (.A(_0519_),
    .ZN(_0520_));
 XNOR2_X1 _4188_ (.A(_0002_),
    .B(_0478_),
    .ZN(_0521_));
 XNOR2_X1 _4189_ (.A(\iir2.y2[7] ),
    .B(_0483_),
    .ZN(_0522_));
 XNOR2_X1 _4190_ (.A(_0519_),
    .B(_0521_),
    .ZN(_0523_));
 INV_X1 _4191_ (.A(_0523_),
    .ZN(_0524_));
 OAI22_X1 _4192_ (.A1(_0520_),
    .A2(_0521_),
    .B1(_0522_),
    .B2(_0524_),
    .ZN(_0525_));
 XNOR2_X1 _4193_ (.A(_0484_),
    .B(_0510_),
    .ZN(_0526_));
 AND2_X1 _4194_ (.A1(_0525_),
    .A2(_0526_),
    .ZN(_0527_));
 INV_X1 _4195_ (.A(_0489_),
    .ZN(_0528_));
 AOI21_X1 _4196_ (.A(_0528_),
    .B1(_0483_),
    .B2(\iir2.y2[7] ),
    .ZN(_0529_));
 XNOR2_X1 _4197_ (.A(\iir2.y2[4] ),
    .B(_0529_),
    .ZN(_0530_));
 XOR2_X1 _4198_ (.A(_0525_),
    .B(_0526_),
    .Z(_0531_));
 AOI21_X1 _4199_ (.A(_0527_),
    .B1(_0530_),
    .B2(_0531_),
    .ZN(_0532_));
 XOR2_X1 _4200_ (.A(_0028_),
    .B(_0489_),
    .Z(_0533_));
 OAI21_X1 _4201_ (.A(_0511_),
    .B1(_0512_),
    .B2(_0452_),
    .ZN(_0534_));
 AOI21_X1 _4202_ (.A(_0533_),
    .B1(_0534_),
    .B2(_0488_),
    .ZN(_0535_));
 OR3_X1 _4203_ (.A1(_0514_),
    .A2(_0532_),
    .A3(_0535_),
    .ZN(_0536_));
 INV_X1 _4204_ (.A(\iir2.y2[4] ),
    .ZN(_0537_));
 OR2_X1 _4205_ (.A1(_0537_),
    .A2(_0529_),
    .ZN(_0538_));
 XNOR2_X1 _4206_ (.A(\iir2.y2[2] ),
    .B(_0538_),
    .ZN(_0539_));
 OAI21_X1 _4207_ (.A(_0490_),
    .B1(_0491_),
    .B2(_0513_),
    .ZN(_0540_));
 NAND3_X1 _4208_ (.A1(_0488_),
    .A2(_0533_),
    .A3(_0534_),
    .ZN(_0541_));
 AOI221_X1 _4209_ (.A(_0527_),
    .B1(_0530_),
    .B2(_0531_),
    .C1(_0540_),
    .C2(_0541_),
    .ZN(_0542_));
 OAI21_X1 _4210_ (.A(_0536_),
    .B1(_0539_),
    .B2(_0542_),
    .ZN(_0543_));
 OAI21_X1 _4211_ (.A(_0498_),
    .B1(_0499_),
    .B2(_0494_),
    .ZN(_0544_));
 NAND3_X1 _4212_ (.A1(_0500_),
    .A2(_0543_),
    .A3(_0544_),
    .ZN(_0545_));
 AND3_X1 _4213_ (.A1(_0500_),
    .A2(_0543_),
    .A3(_0544_),
    .ZN(_0546_));
 AOI21_X1 _4214_ (.A(_0543_),
    .B1(_0544_),
    .B2(_0500_),
    .ZN(_0547_));
 OR4_X1 _4215_ (.A1(\iir2.y2[2] ),
    .A2(_0538_),
    .A3(_0546_),
    .A4(_0547_),
    .ZN(_0548_));
 AND2_X1 _4216_ (.A1(_0545_),
    .A2(_0548_),
    .ZN(_0549_));
 XNOR2_X1 _4217_ (.A(_0505_),
    .B(_0504_),
    .ZN(_0550_));
 OR2_X1 _4218_ (.A1(_0549_),
    .A2(_0550_),
    .ZN(_0551_));
 AND2_X1 _4219_ (.A1(_0549_),
    .A2(_0550_),
    .ZN(_0552_));
 NOR3_X1 _4220_ (.A1(_0514_),
    .A2(_0532_),
    .A3(_0535_),
    .ZN(_0553_));
 OR3_X1 _4221_ (.A1(_0553_),
    .A2(_0539_),
    .A3(_0542_),
    .ZN(_0554_));
 XNOR2_X1 _4222_ (.A(_0522_),
    .B(_0523_),
    .ZN(_0555_));
 XOR2_X1 _4223_ (.A(\iir2.y2[7] ),
    .B(\iir2.y2[6] ),
    .Z(_0556_));
 INV_X1 _4224_ (.A(_0556_),
    .ZN(_0557_));
 OAI21_X1 _4225_ (.A(_2896_),
    .B1(_2908_),
    .B2(_2909_),
    .ZN(_0558_));
 XOR2_X1 _4226_ (.A(_2898_),
    .B(_0558_),
    .Z(_0559_));
 OR2_X1 _4227_ (.A1(_0518_),
    .A2(_0559_),
    .ZN(_0560_));
 XNOR2_X1 _4228_ (.A(_0518_),
    .B(_0559_),
    .ZN(_0561_));
 INV_X1 _4229_ (.A(_0561_),
    .ZN(_0562_));
 NAND2_X1 _4230_ (.A1(\iir2.y2[7] ),
    .A2(_0562_),
    .ZN(_0563_));
 NAND2_X1 _4231_ (.A1(_0560_),
    .A2(_0563_),
    .ZN(_0564_));
 XNOR2_X1 _4232_ (.A(_0518_),
    .B(_0517_),
    .ZN(_0565_));
 XOR2_X1 _4233_ (.A(_0564_),
    .B(_0565_),
    .Z(_0566_));
 NOR2_X1 _4234_ (.A1(_0557_),
    .A2(_0566_),
    .ZN(_0567_));
 AOI21_X1 _4235_ (.A(_0565_),
    .B1(_0563_),
    .B2(_0560_),
    .ZN(_0568_));
 OAI21_X1 _4236_ (.A(_0555_),
    .B1(_0567_),
    .B2(_0568_),
    .ZN(_0569_));
 NAND3_X1 _4237_ (.A1(_0560_),
    .A2(_0563_),
    .A3(_0565_),
    .ZN(_0570_));
 AOI21_X1 _4238_ (.A(_0568_),
    .B1(_0556_),
    .B2(_0570_),
    .ZN(_0571_));
 XNOR2_X1 _4239_ (.A(_0571_),
    .B(_0555_),
    .ZN(_0572_));
 NAND3_X1 _4240_ (.A1(\iir2.y2[7] ),
    .A2(\iir2.y2[6] ),
    .A3(_0572_),
    .ZN(_0573_));
 AND2_X1 _4241_ (.A1(_0569_),
    .A2(_0573_),
    .ZN(_0574_));
 XNOR2_X1 _4242_ (.A(_0530_),
    .B(_0531_),
    .ZN(_0575_));
 OR2_X1 _4243_ (.A1(_0574_),
    .A2(_0575_),
    .ZN(_0576_));
 NOR2_X1 _4244_ (.A1(\iir2.y2[1] ),
    .A2(\iir2.y2[0] ),
    .ZN(_0577_));
 NAND2_X1 _4245_ (.A1(\iir2.y2[3] ),
    .A2(_0577_),
    .ZN(_0578_));
 OAI21_X1 _4246_ (.A(\iir2.y2[1] ),
    .B1(\iir2.y2[0] ),
    .B2(_0496_),
    .ZN(_0579_));
 AND2_X1 _4247_ (.A1(_0578_),
    .A2(_0579_),
    .ZN(_0580_));
 INV_X1 _4248_ (.A(_0580_),
    .ZN(_0581_));
 XNOR2_X1 _4249_ (.A(_0574_),
    .B(_0575_),
    .ZN(_0582_));
 OAI21_X1 _4250_ (.A(_0576_),
    .B1(_0581_),
    .B2(_0582_),
    .ZN(_0583_));
 OAI21_X1 _4251_ (.A(_0539_),
    .B1(_0542_),
    .B2(_0553_),
    .ZN(_0584_));
 NAND3_X1 _4252_ (.A1(_0554_),
    .A2(_0583_),
    .A3(_0584_),
    .ZN(_0585_));
 AOI21_X1 _4253_ (.A(_0583_),
    .B1(_0584_),
    .B2(_0554_),
    .ZN(_0586_));
 OAI21_X1 _4254_ (.A(_0585_),
    .B1(_0586_),
    .B2(_0578_),
    .ZN(_0587_));
 OAI22_X1 _4255_ (.A1(\iir2.y2[2] ),
    .A2(_0538_),
    .B1(_0546_),
    .B2(_0547_),
    .ZN(_0588_));
 AND3_X1 _4256_ (.A1(_0548_),
    .A2(_0587_),
    .A3(_0588_),
    .ZN(_0589_));
 AOI21_X1 _4257_ (.A(_0587_),
    .B1(_0588_),
    .B2(_0548_),
    .ZN(_0590_));
 INV_X1 _4258_ (.A(_0590_),
    .ZN(_0591_));
 AND3_X1 _4259_ (.A1(_0554_),
    .A2(_0583_),
    .A3(_0584_),
    .ZN(_0592_));
 OR3_X1 _4260_ (.A1(_0578_),
    .A2(_0592_),
    .A3(_0586_),
    .ZN(_0593_));
 XNOR2_X1 _4261_ (.A(_0556_),
    .B(_0566_),
    .ZN(_0594_));
 XNOR2_X1 _4262_ (.A(\iir2.y2[6] ),
    .B(\iir2.y2[5] ),
    .ZN(_0595_));
 XOR2_X1 _4263_ (.A(_2908_),
    .B(_2909_),
    .Z(_0596_));
 NAND2_X1 _4264_ (.A1(\iir2.y2[7] ),
    .A2(_0596_),
    .ZN(_0597_));
 XNOR2_X1 _4265_ (.A(\iir2.y2[7] ),
    .B(_0596_),
    .ZN(_0598_));
 OAI21_X1 _4266_ (.A(_0597_),
    .B1(_0598_),
    .B2(_0297_),
    .ZN(_0599_));
 INV_X1 _4267_ (.A(_0599_),
    .ZN(_0600_));
 XOR2_X1 _4268_ (.A(\iir2.y2[7] ),
    .B(_0561_),
    .Z(_0601_));
 XNOR2_X1 _4269_ (.A(_0600_),
    .B(_0601_),
    .ZN(_0602_));
 NOR2_X1 _4270_ (.A1(_0595_),
    .A2(_0602_),
    .ZN(_0603_));
 NOR2_X1 _4271_ (.A1(_0600_),
    .A2(_0601_),
    .ZN(_0604_));
 OAI21_X1 _4272_ (.A(_0594_),
    .B1(_0603_),
    .B2(_0604_),
    .ZN(_0605_));
 NAND2_X1 _4273_ (.A1(\iir2.y2[6] ),
    .A2(\iir2.y2[5] ),
    .ZN(_0606_));
 XNOR2_X1 _4274_ (.A(_0025_),
    .B(_0606_),
    .ZN(_0607_));
 NOR2_X1 _4275_ (.A1(_0604_),
    .A2(_0603_),
    .ZN(_0608_));
 XOR2_X1 _4276_ (.A(_0608_),
    .B(_0594_),
    .Z(_0609_));
 OAI21_X1 _4277_ (.A(_0605_),
    .B1(_0607_),
    .B2(_0609_),
    .ZN(_0610_));
 NAND2_X1 _4278_ (.A1(\iir2.y2[7] ),
    .A2(\iir2.y2[6] ),
    .ZN(_0611_));
 XNOR2_X1 _4279_ (.A(_0611_),
    .B(_0572_),
    .ZN(_0612_));
 NAND2_X1 _4280_ (.A1(_0610_),
    .A2(_0612_),
    .ZN(_0613_));
 XOR2_X1 _4281_ (.A(\iir2.y2[3] ),
    .B(\iir2.y2[0] ),
    .Z(_0614_));
 OAI21_X1 _4282_ (.A(_0614_),
    .B1(_0606_),
    .B2(_0025_),
    .ZN(_0615_));
 OR3_X1 _4283_ (.A1(_0025_),
    .A2(_0606_),
    .A3(_0614_),
    .ZN(_0616_));
 NAND2_X1 _4284_ (.A1(_0615_),
    .A2(_0616_),
    .ZN(_0617_));
 XNOR2_X1 _4285_ (.A(_0610_),
    .B(_0612_),
    .ZN(_0618_));
 OAI21_X1 _4286_ (.A(_0613_),
    .B1(_0617_),
    .B2(_0618_),
    .ZN(_0619_));
 XNOR2_X1 _4287_ (.A(_0580_),
    .B(_0582_),
    .ZN(_0620_));
 NAND2_X1 _4288_ (.A1(_0619_),
    .A2(_0620_),
    .ZN(_0621_));
 XNOR2_X1 _4289_ (.A(_0619_),
    .B(_0620_),
    .ZN(_0622_));
 OAI21_X1 _4290_ (.A(_0621_),
    .B1(_0622_),
    .B2(_0616_),
    .ZN(_0623_));
 OAI21_X1 _4291_ (.A(_0578_),
    .B1(_0592_),
    .B2(_0586_),
    .ZN(_0624_));
 AND3_X1 _4292_ (.A1(_0593_),
    .A2(_0623_),
    .A3(_0624_),
    .ZN(_0625_));
 NAND2_X1 _4293_ (.A1(\iir2.y2[5] ),
    .A2(\iir2.y2[4] ),
    .ZN(_0626_));
 XOR2_X1 _4294_ (.A(_0027_),
    .B(_0626_),
    .Z(_0627_));
 XNOR2_X1 _4295_ (.A(_2906_),
    .B(_2907_),
    .ZN(_0628_));
 XNOR2_X1 _4296_ (.A(_0297_),
    .B(_0628_),
    .ZN(_0629_));
 OAI22_X1 _4297_ (.A1(_0026_),
    .A2(_0628_),
    .B1(_0629_),
    .B2(_0426_),
    .ZN(_0630_));
 XNOR2_X1 _4298_ (.A(_0297_),
    .B(_0598_),
    .ZN(_0631_));
 INV_X1 _4299_ (.A(_0631_),
    .ZN(_0632_));
 NAND2_X1 _4300_ (.A1(_0630_),
    .A2(_0632_),
    .ZN(_0633_));
 XNOR2_X1 _4301_ (.A(\iir2.y2[5] ),
    .B(\iir2.y2[4] ),
    .ZN(_0634_));
 XOR2_X1 _4302_ (.A(_0630_),
    .B(_0631_),
    .Z(_0635_));
 OAI21_X1 _4303_ (.A(_0633_),
    .B1(_0634_),
    .B2(_0635_),
    .ZN(_0636_));
 XOR2_X1 _4304_ (.A(_0595_),
    .B(_0602_),
    .Z(_0637_));
 XOR2_X1 _4305_ (.A(_0636_),
    .B(_0637_),
    .Z(_0638_));
 AND2_X1 _4306_ (.A1(_0627_),
    .A2(_0638_),
    .ZN(_0639_));
 AOI21_X1 _4307_ (.A(_0639_),
    .B1(_0637_),
    .B2(_0636_),
    .ZN(_0640_));
 XNOR2_X1 _4308_ (.A(_0607_),
    .B(_0609_),
    .ZN(_0641_));
 OR2_X1 _4309_ (.A1(_0640_),
    .A2(_0641_),
    .ZN(_0642_));
 INV_X1 _4310_ (.A(_0642_),
    .ZN(_0643_));
 XNOR2_X1 _4311_ (.A(_0640_),
    .B(_0641_),
    .ZN(_0644_));
 NOR3_X1 _4312_ (.A1(_0027_),
    .A2(_0626_),
    .A3(_0644_),
    .ZN(_0645_));
 NOR2_X1 _4313_ (.A1(_0643_),
    .A2(_0645_),
    .ZN(_0646_));
 XNOR2_X1 _4314_ (.A(_0617_),
    .B(_0618_),
    .ZN(_0647_));
 OR2_X1 _4315_ (.A1(_0646_),
    .A2(_0647_),
    .ZN(_0648_));
 INV_X1 _4316_ (.A(_0648_),
    .ZN(_0649_));
 XOR2_X1 _4317_ (.A(_0616_),
    .B(_0622_),
    .Z(_0650_));
 NAND2_X1 _4318_ (.A1(_0649_),
    .A2(_0650_),
    .ZN(_0651_));
 XNOR2_X1 _4319_ (.A(_0649_),
    .B(_0650_),
    .ZN(_0652_));
 NOR2_X1 _4320_ (.A1(_0027_),
    .A2(_0626_),
    .ZN(_0653_));
 XNOR2_X1 _4321_ (.A(_0653_),
    .B(_0644_),
    .ZN(_0654_));
 NAND2_X1 _4322_ (.A1(\iir2.y2[4] ),
    .A2(\iir2.y2[3] ),
    .ZN(_0655_));
 NOR2_X1 _4323_ (.A1(_0029_),
    .A2(_0655_),
    .ZN(_0656_));
 XNOR2_X1 _4324_ (.A(_0627_),
    .B(_0638_),
    .ZN(_0657_));
 XOR2_X1 _4325_ (.A(_0029_),
    .B(_0655_),
    .Z(_0658_));
 XNOR2_X1 _4326_ (.A(_2904_),
    .B(_2905_),
    .ZN(_0659_));
 XNOR2_X1 _4327_ (.A(_0426_),
    .B(_0659_),
    .ZN(_0660_));
 OAI22_X1 _4328_ (.A1(_0028_),
    .A2(_0659_),
    .B1(_0660_),
    .B2(_0537_),
    .ZN(_0661_));
 XNOR2_X1 _4329_ (.A(\iir2.y2[5] ),
    .B(_0629_),
    .ZN(_0662_));
 NAND2_X1 _4330_ (.A1(_0661_),
    .A2(_0662_),
    .ZN(_0663_));
 XNOR2_X1 _4331_ (.A(\iir2.y2[4] ),
    .B(\iir2.y2[3] ),
    .ZN(_0664_));
 XNOR2_X1 _4332_ (.A(_0661_),
    .B(_0662_),
    .ZN(_0665_));
 OAI21_X1 _4333_ (.A(_0663_),
    .B1(_0664_),
    .B2(_0665_),
    .ZN(_0666_));
 XOR2_X1 _4334_ (.A(_0634_),
    .B(_0635_),
    .Z(_0667_));
 XNOR2_X1 _4335_ (.A(_0666_),
    .B(_0667_),
    .ZN(_0668_));
 INV_X1 _4336_ (.A(_0668_),
    .ZN(_0669_));
 NAND2_X1 _4337_ (.A1(_0658_),
    .A2(_0669_),
    .ZN(_0670_));
 NAND2_X1 _4338_ (.A1(_0666_),
    .A2(_0667_),
    .ZN(_0671_));
 AOI21_X1 _4339_ (.A(_0657_),
    .B1(_0670_),
    .B2(_0671_),
    .ZN(_0672_));
 AND3_X1 _4340_ (.A1(_0671_),
    .A2(_0670_),
    .A3(_0657_),
    .ZN(_0673_));
 NOR2_X1 _4341_ (.A1(_0672_),
    .A2(_0673_),
    .ZN(_0674_));
 AND2_X1 _4342_ (.A1(_0656_),
    .A2(_0674_),
    .ZN(_0675_));
 OAI21_X1 _4343_ (.A(_0654_),
    .B1(_0675_),
    .B2(_0672_),
    .ZN(_0676_));
 XNOR2_X1 _4344_ (.A(_0646_),
    .B(_0647_),
    .ZN(_0677_));
 NOR2_X1 _4345_ (.A1(_0676_),
    .A2(_0677_),
    .ZN(_0678_));
 OR3_X1 _4346_ (.A1(_0672_),
    .A2(_0675_),
    .A3(_0654_),
    .ZN(_0679_));
 NAND2_X1 _4347_ (.A1(_0676_),
    .A2(_0679_),
    .ZN(_0680_));
 XOR2_X1 _4348_ (.A(_0664_),
    .B(_0665_),
    .Z(_0681_));
 XNOR2_X1 _4349_ (.A(\iir2.y2[3] ),
    .B(\iir2.y2[2] ),
    .ZN(_0682_));
 XOR2_X1 _4350_ (.A(_2902_),
    .B(_2903_),
    .Z(_0683_));
 NAND2_X1 _4351_ (.A1(\iir2.y2[4] ),
    .A2(_0683_),
    .ZN(_0684_));
 XNOR2_X1 _4352_ (.A(\iir2.y2[4] ),
    .B(_0683_),
    .ZN(_0685_));
 OAI21_X1 _4353_ (.A(_0684_),
    .B1(_0685_),
    .B2(_0496_),
    .ZN(_0686_));
 XNOR2_X1 _4354_ (.A(\iir2.y2[4] ),
    .B(_0660_),
    .ZN(_0687_));
 XNOR2_X1 _4355_ (.A(_0686_),
    .B(_0687_),
    .ZN(_0688_));
 NOR2_X1 _4356_ (.A1(_0682_),
    .A2(_0688_),
    .ZN(_0689_));
 AND2_X1 _4357_ (.A1(_0686_),
    .A2(_0687_),
    .ZN(_0690_));
 OAI21_X1 _4358_ (.A(_0681_),
    .B1(_0689_),
    .B2(_0690_),
    .ZN(_0691_));
 OR3_X1 _4359_ (.A1(_0690_),
    .A2(_0689_),
    .A3(_0681_),
    .ZN(_0692_));
 NAND2_X1 _4360_ (.A1(_0691_),
    .A2(_0692_),
    .ZN(_0693_));
 NAND2_X1 _4361_ (.A1(\iir2.y2[3] ),
    .A2(\iir2.y2[2] ),
    .ZN(_0694_));
 OAI21_X1 _4362_ (.A(_0691_),
    .B1(_0693_),
    .B2(_0694_),
    .ZN(_0695_));
 XNOR2_X1 _4363_ (.A(_0658_),
    .B(_0668_),
    .ZN(_0696_));
 XOR2_X1 _4364_ (.A(_0656_),
    .B(_0674_),
    .Z(_0697_));
 NAND3_X1 _4365_ (.A1(_0695_),
    .A2(_0696_),
    .A3(_0697_),
    .ZN(_0698_));
 XNOR2_X1 _4366_ (.A(_2849_),
    .B(_2901_),
    .ZN(_0699_));
 NOR2_X1 _4367_ (.A1(_0496_),
    .A2(_0699_),
    .ZN(_0700_));
 INV_X1 _4368_ (.A(\iir2.y2[2] ),
    .ZN(_0701_));
 XNOR2_X1 _4369_ (.A(_0496_),
    .B(_0699_),
    .ZN(_0702_));
 NOR2_X1 _4370_ (.A1(_0701_),
    .A2(_0702_),
    .ZN(_0703_));
 NOR2_X1 _4371_ (.A1(_0700_),
    .A2(_0703_),
    .ZN(_0704_));
 XNOR2_X1 _4372_ (.A(_0496_),
    .B(_0685_),
    .ZN(_0705_));
 NOR2_X1 _4373_ (.A1(_0704_),
    .A2(_0705_),
    .ZN(_0706_));
 XOR2_X1 _4374_ (.A(\iir2.y2[2] ),
    .B(\iir2.y2[1] ),
    .Z(_0707_));
 XOR2_X1 _4375_ (.A(_0704_),
    .B(_0705_),
    .Z(_0708_));
 AOI21_X1 _4376_ (.A(_0706_),
    .B1(_0707_),
    .B2(_0708_),
    .ZN(_0709_));
 XNOR2_X1 _4377_ (.A(_0682_),
    .B(_0688_),
    .ZN(_0710_));
 XOR2_X1 _4378_ (.A(_0709_),
    .B(_0710_),
    .Z(_0711_));
 NAND3_X1 _4379_ (.A1(\iir2.y2[2] ),
    .A2(\iir2.y2[1] ),
    .A3(_0711_),
    .ZN(_0712_));
 OAI21_X1 _4380_ (.A(_0712_),
    .B1(_0710_),
    .B2(_0709_),
    .ZN(_0713_));
 XOR2_X1 _4381_ (.A(_0694_),
    .B(_0693_),
    .Z(_0714_));
 NAND2_X1 _4382_ (.A1(_0713_),
    .A2(_0714_),
    .ZN(_0715_));
 NOR2_X1 _4383_ (.A1(_0713_),
    .A2(_0714_),
    .ZN(_0716_));
 AND2_X1 _4384_ (.A1(\iir2.y2[1] ),
    .A2(\iir2.y2[0] ),
    .ZN(_0717_));
 OR2_X1 _4385_ (.A1(_0577_),
    .A2(_0717_),
    .ZN(_0718_));
 NAND2_X1 _4386_ (.A1(\iir2.x2[0] ),
    .A2(_2401_),
    .ZN(_0719_));
 XOR2_X1 _4387_ (.A(_2393_),
    .B(_0719_),
    .Z(_0720_));
 XNOR2_X1 _4388_ (.A(_0701_),
    .B(_0720_),
    .ZN(_0721_));
 INV_X1 _4389_ (.A(\iir2.y2[1] ),
    .ZN(_0722_));
 OAI22_X1 _4390_ (.A1(_0025_),
    .A2(_0720_),
    .B1(_0721_),
    .B2(_0722_),
    .ZN(_0723_));
 XNOR2_X1 _4391_ (.A(\iir2.y2[2] ),
    .B(_0702_),
    .ZN(_0724_));
 XNOR2_X1 _4392_ (.A(_0723_),
    .B(_0724_),
    .ZN(_0725_));
 NOR2_X1 _4393_ (.A1(_0718_),
    .A2(_0725_),
    .ZN(_0726_));
 AOI21_X1 _4394_ (.A(_0726_),
    .B1(_0724_),
    .B2(_0723_),
    .ZN(_0727_));
 XNOR2_X1 _4395_ (.A(_0707_),
    .B(_0708_),
    .ZN(_0728_));
 NOR2_X1 _4396_ (.A1(_0727_),
    .A2(_0728_),
    .ZN(_0729_));
 XOR2_X1 _4397_ (.A(_0727_),
    .B(_0728_),
    .Z(_0730_));
 AOI21_X1 _4398_ (.A(_0729_),
    .B1(_0730_),
    .B2(_0717_),
    .ZN(_0731_));
 NAND2_X1 _4399_ (.A1(\iir2.y2[2] ),
    .A2(\iir2.y2[1] ),
    .ZN(_0732_));
 XOR2_X1 _4400_ (.A(_0732_),
    .B(_0711_),
    .Z(_0733_));
 NOR2_X1 _4401_ (.A1(_0731_),
    .A2(_0733_),
    .ZN(_0734_));
 NAND2_X1 _4402_ (.A1(_0731_),
    .A2(_0733_),
    .ZN(_0735_));
 NOR2_X1 _4403_ (.A1(_0717_),
    .A2(_0730_),
    .ZN(_0736_));
 INV_X1 _4404_ (.A(\iir1.y[0] ),
    .ZN(_0737_));
 NAND2_X1 _4405_ (.A1(_0737_),
    .A2(\iir2.x2[0] ),
    .ZN(_0738_));
 XNOR2_X1 _4406_ (.A(_2388_),
    .B(_0738_),
    .ZN(_0739_));
 XNOR2_X1 _4407_ (.A(\iir2.y2[1] ),
    .B(_0739_),
    .ZN(_0740_));
 NAND2_X1 _4408_ (.A1(\iir2.y2[0] ),
    .A2(_0740_),
    .ZN(_0741_));
 OAI21_X1 _4409_ (.A(_0741_),
    .B1(_0739_),
    .B2(_0027_),
    .ZN(_0742_));
 INV_X1 _4410_ (.A(_0742_),
    .ZN(_0743_));
 XNOR2_X1 _4411_ (.A(_0722_),
    .B(_0721_),
    .ZN(_0744_));
 NOR2_X1 _4412_ (.A1(_0743_),
    .A2(_0744_),
    .ZN(_0745_));
 XNOR2_X1 _4413_ (.A(\iir1.y[0] ),
    .B(\iir2.x2[0] ),
    .ZN(_0746_));
 XNOR2_X1 _4414_ (.A(\iir2.y2[0] ),
    .B(_0740_),
    .ZN(_0747_));
 XNOR2_X1 _4415_ (.A(_0742_),
    .B(_0744_),
    .ZN(_0748_));
 XNOR2_X1 _4416_ (.A(\iir2.y2[0] ),
    .B(_0748_),
    .ZN(_0749_));
 NOR4_X1 _4417_ (.A1(_0029_),
    .A2(_0746_),
    .A3(_0747_),
    .A4(_0749_),
    .ZN(_0750_));
 NAND2_X1 _4418_ (.A1(_0745_),
    .A2(_0750_),
    .ZN(_0751_));
 AND2_X1 _4419_ (.A1(_0718_),
    .A2(_0725_),
    .ZN(_0752_));
 OAI21_X1 _4420_ (.A(_0751_),
    .B1(_0752_),
    .B2(_0726_),
    .ZN(_0753_));
 NAND2_X1 _4421_ (.A1(\iir2.y2[0] ),
    .A2(_0748_),
    .ZN(_0754_));
 OAI21_X1 _4422_ (.A(_0754_),
    .B1(_0744_),
    .B2(_0743_),
    .ZN(_0755_));
 OAI21_X1 _4423_ (.A(_0753_),
    .B1(_0755_),
    .B2(_0750_),
    .ZN(_0756_));
 AOI211_X1 _4424_ (.A(_0736_),
    .B(_0756_),
    .C1(_0717_),
    .C2(_0730_),
    .ZN(_0757_));
 AOI21_X1 _4425_ (.A(_0734_),
    .B1(_0735_),
    .B2(_0757_),
    .ZN(_0758_));
 OAI21_X1 _4426_ (.A(_0715_),
    .B1(_0716_),
    .B2(_0758_),
    .ZN(_0759_));
 NAND2_X1 _4427_ (.A1(_0695_),
    .A2(_0696_),
    .ZN(_0760_));
 OR2_X1 _4428_ (.A1(_0695_),
    .A2(_0696_),
    .ZN(_0761_));
 NAND4_X1 _4429_ (.A1(_0759_),
    .A2(_0760_),
    .A3(_0697_),
    .A4(_0761_),
    .ZN(_0762_));
 AOI21_X1 _4430_ (.A(_0680_),
    .B1(_0698_),
    .B2(_0762_),
    .ZN(_0763_));
 XOR2_X1 _4431_ (.A(_0676_),
    .B(_0677_),
    .Z(_0764_));
 AOI21_X1 _4432_ (.A(_0678_),
    .B1(_0763_),
    .B2(_0764_),
    .ZN(_0765_));
 OAI21_X1 _4433_ (.A(_0651_),
    .B1(_0652_),
    .B2(_0765_),
    .ZN(_0766_));
 AOI21_X1 _4434_ (.A(_0623_),
    .B1(_0624_),
    .B2(_0593_),
    .ZN(_0767_));
 NOR4_X1 _4435_ (.A1(_0589_),
    .A2(_0590_),
    .A3(_0625_),
    .A4(_0767_),
    .ZN(_0768_));
 AOI221_X1 _4436_ (.A(_0589_),
    .B1(_0591_),
    .B2(_0625_),
    .C1(_0766_),
    .C2(_0768_),
    .ZN(_0769_));
 OAI21_X1 _4437_ (.A(_0551_),
    .B1(_0552_),
    .B2(_0769_),
    .ZN(_0770_));
 AOI21_X1 _4438_ (.A(_0508_),
    .B1(_0509_),
    .B2(_0770_),
    .ZN(_0771_));
 OAI21_X1 _4439_ (.A(_0475_),
    .B1(_0477_),
    .B2(_0771_),
    .ZN(_0772_));
 XNOR2_X1 _4440_ (.A(_0364_),
    .B(_0415_),
    .ZN(_0773_));
 AOI21_X1 _4441_ (.A(_0416_),
    .B1(_0772_),
    .B2(_0773_),
    .ZN(_0774_));
 NAND2_X1 _4442_ (.A1(_0366_),
    .A2(_0414_),
    .ZN(_0775_));
 OAI21_X1 _4443_ (.A(_0775_),
    .B1(_0413_),
    .B2(_0368_),
    .ZN(_0776_));
 NOR2_X1 _4444_ (.A1(_0440_),
    .A2(\iir2.y2[8] ),
    .ZN(_0777_));
 INV_X1 _4445_ (.A(_0357_),
    .ZN(_0778_));
 NAND2_X1 _4446_ (.A1(_0293_),
    .A2(_0778_),
    .ZN(_0779_));
 NOR3_X1 _4447_ (.A1(_0002_),
    .A2(_0411_),
    .A3(_0779_),
    .ZN(_0780_));
 AND2_X1 _4448_ (.A1(_1308_),
    .A2(_0412_),
    .ZN(_0781_));
 NOR2_X1 _4449_ (.A1(_0780_),
    .A2(_0781_),
    .ZN(_0782_));
 NOR3_X1 _4450_ (.A1(_0002_),
    .A2(_0778_),
    .A3(_0411_),
    .ZN(_0783_));
 OAI21_X1 _4451_ (.A(_0440_),
    .B1(_0408_),
    .B2(_0409_),
    .ZN(_0784_));
 OR3_X1 _4452_ (.A1(_0440_),
    .A2(_0408_),
    .A3(_0409_),
    .ZN(_0785_));
 AOI21_X1 _4453_ (.A(_0002_),
    .B1(_0784_),
    .B2(_0785_),
    .ZN(_0786_));
 NOR2_X1 _4454_ (.A1(_0347_),
    .A2(_0405_),
    .ZN(_0787_));
 AOI21_X1 _4455_ (.A(_0787_),
    .B1(_0406_),
    .B2(_0370_),
    .ZN(_0788_));
 NAND3_X1 _4456_ (.A1(_0349_),
    .A2(_0353_),
    .A3(_0406_),
    .ZN(_0789_));
 NOR2_X1 _4457_ (.A1(_2845_),
    .A2(_0225_),
    .ZN(_0790_));
 AOI21_X1 _4458_ (.A(_0227_),
    .B1(_0790_),
    .B2(_0220_),
    .ZN(_0791_));
 NAND4_X1 _4459_ (.A1(_0214_),
    .A2(_0291_),
    .A3(_0349_),
    .A4(_0406_),
    .ZN(_0792_));
 OR2_X1 _4460_ (.A1(_0791_),
    .A2(_0792_),
    .ZN(_0793_));
 NOR3_X1 _4461_ (.A1(_2864_),
    .A2(_2866_),
    .A3(_2916_),
    .ZN(_0794_));
 NAND2_X1 _4462_ (.A1(_0794_),
    .A2(_0790_),
    .ZN(_0795_));
 OR3_X1 _4463_ (.A1(_2913_),
    .A2(_0795_),
    .A3(_0792_),
    .ZN(_0796_));
 AND4_X1 _4464_ (.A1(_0788_),
    .A2(_0789_),
    .A3(_0793_),
    .A4(_0796_),
    .ZN(_0797_));
 AOI21_X1 _4465_ (.A(_0404_),
    .B1(_0373_),
    .B2(_0372_),
    .ZN(_0798_));
 OR3_X1 _4466_ (.A1(z[8]),
    .A2(_0251_),
    .A3(_0403_),
    .ZN(_0799_));
 INV_X1 _4467_ (.A(_0402_),
    .ZN(_0800_));
 OAI21_X1 _4468_ (.A(_0799_),
    .B1(_0800_),
    .B2(_0377_),
    .ZN(_0801_));
 NOR2_X1 _4469_ (.A1(z[9]),
    .A2(_0315_),
    .ZN(_0802_));
 NAND2_X1 _4470_ (.A1(_0379_),
    .A2(_0401_),
    .ZN(_0803_));
 NAND2_X1 _4471_ (.A1(z[10]),
    .A2(_0400_),
    .ZN(_0804_));
 INV_X1 _4472_ (.A(_0804_),
    .ZN(_0805_));
 NAND2_X1 _4473_ (.A1(_0341_),
    .A2(_0805_),
    .ZN(_0806_));
 OAI21_X1 _4474_ (.A(_0803_),
    .B1(_0806_),
    .B2(_0318_),
    .ZN(_0807_));
 NOR2_X1 _4475_ (.A1(_2753_),
    .A2(z[8]),
    .ZN(_0808_));
 XNOR2_X1 _4476_ (.A(_2786_),
    .B(_0808_),
    .ZN(_0809_));
 INV_X1 _4477_ (.A(_0399_),
    .ZN(_0810_));
 NOR2_X1 _4478_ (.A1(_0381_),
    .A2(_0810_),
    .ZN(_0811_));
 AOI21_X1 _4479_ (.A(_0811_),
    .B1(_0398_),
    .B2(_0383_),
    .ZN(_0812_));
 MUX2_X1 _4480_ (.A(_0031_),
    .B(_0385_),
    .S(_0392_),
    .Z(_0813_));
 MUX2_X1 _4481_ (.A(_0394_),
    .B(_0396_),
    .S(_2554_),
    .Z(_0814_));
 XNOR2_X1 _4482_ (.A(_0813_),
    .B(_0814_),
    .ZN(_0815_));
 XNOR2_X1 _4483_ (.A(_0812_),
    .B(_0815_),
    .ZN(_0816_));
 AOI21_X1 _4484_ (.A(_0816_),
    .B1(_0805_),
    .B2(_0341_),
    .ZN(_0817_));
 XNOR2_X1 _4485_ (.A(_0809_),
    .B(_0817_),
    .ZN(_0818_));
 XNOR2_X1 _4486_ (.A(_0807_),
    .B(_0818_),
    .ZN(_0819_));
 XNOR2_X1 _4487_ (.A(_0802_),
    .B(_0819_),
    .ZN(_0820_));
 XOR2_X1 _4488_ (.A(_0801_),
    .B(_0820_),
    .Z(_0821_));
 XNOR2_X1 _4489_ (.A(_0798_),
    .B(_0821_),
    .ZN(_0822_));
 XOR2_X1 _4490_ (.A(_0797_),
    .B(_0822_),
    .Z(_0823_));
 XNOR2_X1 _4491_ (.A(\iir2.y2[10] ),
    .B(_0823_),
    .ZN(_0824_));
 XNOR2_X1 _4492_ (.A(_0786_),
    .B(_0824_),
    .ZN(_0825_));
 XNOR2_X1 _4493_ (.A(_0783_),
    .B(_0825_),
    .ZN(_0826_));
 XNOR2_X1 _4494_ (.A(_0447_),
    .B(_0826_),
    .ZN(_0827_));
 XNOR2_X1 _4495_ (.A(_0782_),
    .B(_0827_),
    .ZN(_0828_));
 XOR2_X1 _4496_ (.A(_0777_),
    .B(_0828_),
    .Z(_0829_));
 XNOR2_X1 _4497_ (.A(_0776_),
    .B(_0829_),
    .ZN(_0830_));
 XOR2_X1 _4498_ (.A(_0774_),
    .B(_0830_),
    .Z(_0831_));
 INV_X1 _4499_ (.A(_0773_),
    .ZN(_0832_));
 XNOR2_X1 _4500_ (.A(_0772_),
    .B(_0832_),
    .ZN(_0833_));
 OR2_X1 _4501_ (.A1(_0472_),
    .A2(_0473_),
    .ZN(_0834_));
 INV_X1 _4502_ (.A(_0476_),
    .ZN(_0835_));
 OAI21_X1 _4503_ (.A(_0834_),
    .B1(_0771_),
    .B2(_0835_),
    .ZN(_0836_));
 XOR2_X1 _4504_ (.A(_0439_),
    .B(_0836_),
    .Z(_0837_));
 XNOR2_X1 _4505_ (.A(_0771_),
    .B(_0476_),
    .ZN(_0838_));
 XOR2_X1 _4506_ (.A(_0509_),
    .B(_0770_),
    .Z(_0839_));
 XOR2_X1 _4507_ (.A(_0549_),
    .B(_0550_),
    .Z(_0840_));
 XNOR2_X1 _4508_ (.A(_0840_),
    .B(_0769_),
    .ZN(_0841_));
 NOR2_X1 _4509_ (.A1(_0625_),
    .A2(_0767_),
    .ZN(_0842_));
 XOR2_X1 _4510_ (.A(_0842_),
    .B(_0766_),
    .Z(_0843_));
 NAND3_X1 _4511_ (.A1(_0680_),
    .A2(_0698_),
    .A3(_0762_),
    .ZN(_0844_));
 NAND2_X1 _4512_ (.A1(_0764_),
    .A2(_0844_),
    .ZN(_0845_));
 NOR2_X1 _4513_ (.A1(_0763_),
    .A2(_0845_),
    .ZN(_0846_));
 XOR2_X1 _4514_ (.A(_0652_),
    .B(_0765_),
    .Z(_0847_));
 AND2_X1 _4515_ (.A1(_0846_),
    .A2(_0847_),
    .ZN(_0848_));
 AND2_X1 _4516_ (.A1(_0843_),
    .A2(_0848_),
    .ZN(_0849_));
 OR2_X1 _4517_ (.A1(_0589_),
    .A2(_0590_),
    .ZN(_0850_));
 AOI21_X1 _4518_ (.A(_0625_),
    .B1(_0842_),
    .B2(_0766_),
    .ZN(_0851_));
 XOR2_X1 _4519_ (.A(_0850_),
    .B(_0851_),
    .Z(_0852_));
 AND2_X1 _4520_ (.A1(_0849_),
    .A2(_0852_),
    .ZN(_0853_));
 AND2_X1 _4521_ (.A1(_0841_),
    .A2(_0853_),
    .ZN(_0854_));
 AND2_X1 _4522_ (.A1(_0839_),
    .A2(_0854_),
    .ZN(_0855_));
 AND4_X1 _4523_ (.A1(_0833_),
    .A2(_0837_),
    .A3(_0838_),
    .A4(_0855_),
    .ZN(_0856_));
 OAI21_X1 _4524_ (.A(_1297_),
    .B1(_0831_),
    .B2(_0856_),
    .ZN(_0857_));
 AOI21_X1 _4525_ (.A(_0857_),
    .B1(_0856_),
    .B2(_0831_),
    .ZN(_0119_));
 AND2_X1 _4526_ (.A1(_0838_),
    .A2(_0855_),
    .ZN(_0858_));
 AOI21_X1 _4527_ (.A(_0833_),
    .B1(_0837_),
    .B2(_0858_),
    .ZN(_0859_));
 NOR3_X1 _4528_ (.A1(rst),
    .A2(_0856_),
    .A3(_0859_),
    .ZN(_0118_));
 OAI21_X1 _4529_ (.A(_1297_),
    .B1(_0837_),
    .B2(_0858_),
    .ZN(_0860_));
 AOI21_X1 _4530_ (.A(_0860_),
    .B1(_0858_),
    .B2(_0837_),
    .ZN(_0117_));
 NOR2_X1 _4531_ (.A1(_0838_),
    .A2(_0855_),
    .ZN(_0861_));
 NOR3_X1 _4532_ (.A1(rst),
    .A2(_0858_),
    .A3(_0861_),
    .ZN(_0116_));
 NOR2_X1 _4533_ (.A1(_0839_),
    .A2(_0854_),
    .ZN(_0862_));
 NOR3_X1 _4534_ (.A1(rst),
    .A2(_0855_),
    .A3(_0862_),
    .ZN(_0115_));
 NOR2_X1 _4535_ (.A1(_0841_),
    .A2(_0853_),
    .ZN(_0863_));
 NOR3_X1 _4536_ (.A1(rst),
    .A2(_0854_),
    .A3(_0863_),
    .ZN(_0114_));
 NOR2_X1 _4537_ (.A1(_0849_),
    .A2(_0852_),
    .ZN(_0864_));
 NOR3_X1 _4538_ (.A1(rst),
    .A2(_0853_),
    .A3(_0864_),
    .ZN(_0113_));
 NOR2_X1 _4539_ (.A1(_0843_),
    .A2(_0848_),
    .ZN(_0865_));
 NOR3_X1 _4540_ (.A1(rst),
    .A2(_0849_),
    .A3(_0865_),
    .ZN(_0112_));
 NOR2_X1 _4541_ (.A1(_0846_),
    .A2(_0847_),
    .ZN(_0866_));
 NOR3_X1 _4542_ (.A1(rst),
    .A2(_0848_),
    .A3(_0866_),
    .ZN(_0111_));
 NAND2_X1 _4543_ (.A1(_0776_),
    .A2(_0829_),
    .ZN(_0867_));
 NAND2_X1 _4544_ (.A1(_0365_),
    .A2(_0415_),
    .ZN(_0868_));
 OR2_X1 _4545_ (.A1(_0832_),
    .A2(_0830_),
    .ZN(_0869_));
 OAI221_X1 _4546_ (.A(_0867_),
    .B1(_0830_),
    .B2(_0868_),
    .C1(_0869_),
    .C2(_0475_),
    .ZN(_0870_));
 NOR3_X1 _4547_ (.A1(_0771_),
    .A2(_0477_),
    .A3(_0869_),
    .ZN(_0871_));
 NOR2_X1 _4548_ (.A1(_0870_),
    .A2(_0871_),
    .ZN(_0872_));
 OAI21_X1 _4549_ (.A(_0827_),
    .B1(_0781_),
    .B2(_0780_),
    .ZN(_0873_));
 INV_X1 _4550_ (.A(_0873_),
    .ZN(_0874_));
 AOI21_X1 _4551_ (.A(_0874_),
    .B1(_0828_),
    .B2(_0777_),
    .ZN(_0875_));
 NAND2_X1 _4552_ (.A1(_0783_),
    .A2(_0825_),
    .ZN(_0876_));
 OAI21_X1 _4553_ (.A(_0876_),
    .B1(_0826_),
    .B2(_0237_),
    .ZN(_0877_));
 NOR2_X1 _4554_ (.A1(_0797_),
    .A2(_0822_),
    .ZN(_0878_));
 AOI21_X1 _4555_ (.A(_0878_),
    .B1(_0821_),
    .B2(_0798_),
    .ZN(_0879_));
 NAND2_X1 _4556_ (.A1(_0801_),
    .A2(_0820_),
    .ZN(_0880_));
 NOR3_X1 _4557_ (.A1(z[9]),
    .A2(_0315_),
    .A3(_0819_),
    .ZN(_0881_));
 AOI21_X1 _4558_ (.A(_0881_),
    .B1(_0818_),
    .B2(_0807_),
    .ZN(_0882_));
 NOR3_X1 _4559_ (.A1(_0341_),
    .A2(_0804_),
    .A3(_0816_),
    .ZN(_0883_));
 OR2_X1 _4560_ (.A1(_0805_),
    .A2(_0816_),
    .ZN(_0884_));
 AOI21_X1 _4561_ (.A(_0883_),
    .B1(_0884_),
    .B2(_0809_),
    .ZN(_0885_));
 OAI21_X1 _4562_ (.A(z[9]),
    .B1(z[8]),
    .B2(z[10]),
    .ZN(_0886_));
 XNOR2_X1 _4563_ (.A(_0884_),
    .B(_0886_),
    .ZN(_0887_));
 XNOR2_X1 _4564_ (.A(_0885_),
    .B(_0887_),
    .ZN(_0888_));
 XNOR2_X1 _4565_ (.A(_0882_),
    .B(_0888_),
    .ZN(_0889_));
 XNOR2_X1 _4566_ (.A(_0880_),
    .B(_0889_),
    .ZN(_0890_));
 XNOR2_X1 _4567_ (.A(_0879_),
    .B(_0890_),
    .ZN(_0891_));
 NOR2_X1 _4568_ (.A1(_0448_),
    .A2(\iir2.y2[10] ),
    .ZN(_0892_));
 AOI21_X1 _4569_ (.A(_0892_),
    .B1(_0823_),
    .B2(_0448_),
    .ZN(_0893_));
 XNOR2_X1 _4570_ (.A(_0891_),
    .B(_0893_),
    .ZN(_0894_));
 NOR2_X1 _4571_ (.A1(_0440_),
    .A2(\iir2.y2[9] ),
    .ZN(_0895_));
 AOI211_X1 _4572_ (.A(_0002_),
    .B(_0824_),
    .C1(_0785_),
    .C2(_0784_),
    .ZN(_0896_));
 XNOR2_X1 _4573_ (.A(_0895_),
    .B(_0896_),
    .ZN(_0897_));
 XNOR2_X1 _4574_ (.A(_0894_),
    .B(_0897_),
    .ZN(_0898_));
 XOR2_X1 _4575_ (.A(_0877_),
    .B(_0898_),
    .Z(_0899_));
 XNOR2_X1 _4576_ (.A(_0875_),
    .B(_0899_),
    .ZN(_0900_));
 XNOR2_X1 _4577_ (.A(_0872_),
    .B(_0900_),
    .ZN(_0901_));
 AOI21_X1 _4578_ (.A(_0901_),
    .B1(_0856_),
    .B2(_0831_),
    .ZN(_0902_));
 AND3_X1 _4579_ (.A1(_0831_),
    .A2(_0856_),
    .A3(_0901_),
    .ZN(_0903_));
 NOR3_X1 _4580_ (.A1(rst),
    .A2(_0902_),
    .A3(_0903_),
    .ZN(_0110_));
 OR2_X1 _4581_ (.A1(_0764_),
    .A2(_0844_),
    .ZN(_0904_));
 AND3_X1 _4582_ (.A1(_1297_),
    .A2(_0845_),
    .A3(_0904_),
    .ZN(_0109_));
 NOR2_X1 _4583_ (.A1(rst),
    .A2(net64),
    .ZN(_0108_));
 NOR2_X1 _4584_ (.A1(rst),
    .A2(_2613_),
    .ZN(_0107_));
 AND2_X1 _4585_ (.A1(_1297_),
    .A2(net67),
    .ZN(_0106_));
 AND2_X1 _4586_ (.A1(_1297_),
    .A2(net80),
    .ZN(_0105_));
 AND2_X1 _4587_ (.A1(_1297_),
    .A2(net57),
    .ZN(_0104_));
 AND2_X1 _4588_ (.A1(_1297_),
    .A2(net69),
    .ZN(_0103_));
 AND2_X1 _4589_ (.A1(_1297_),
    .A2(net55),
    .ZN(_0102_));
 AND2_X1 _4590_ (.A1(_1297_),
    .A2(net65),
    .ZN(_0101_));
 AND2_X1 _4591_ (.A1(_1297_),
    .A2(net53),
    .ZN(_0100_));
 NOR2_X1 _4592_ (.A1(rst),
    .A2(_2786_),
    .ZN(_0099_));
 NOR2_X1 _4593_ (.A1(rst),
    .A2(net50),
    .ZN(_0098_));
 NOR2_X1 _4594_ (.A1(rst),
    .A2(_2561_),
    .ZN(_0097_));
 NOR2_X1 _4595_ (.A1(rst),
    .A2(net71),
    .ZN(_0096_));
 NOR2_X1 _4596_ (.A1(rst),
    .A2(_2432_),
    .ZN(_0095_));
 NOR2_X1 _4597_ (.A1(rst),
    .A2(net62),
    .ZN(_0094_));
 INV_X1 _4598_ (.A(net88),
    .ZN(_0905_));
 NOR2_X1 _4599_ (.A1(rst),
    .A2(_0905_),
    .ZN(_0093_));
 NOR2_X1 _4600_ (.A1(rst),
    .A2(_2429_),
    .ZN(_0092_));
 INV_X1 _4601_ (.A(net72),
    .ZN(_0906_));
 NOR2_X1 _4602_ (.A1(rst),
    .A2(net73),
    .ZN(_0091_));
 NOR2_X1 _4603_ (.A1(rst),
    .A2(net77),
    .ZN(_0090_));
 NOR2_X1 _4604_ (.A1(rst),
    .A2(_1407_),
    .ZN(_0089_));
 NOR2_X1 _4605_ (.A1(rst),
    .A2(_2704_),
    .ZN(_0088_));
 NOR2_X1 _4606_ (.A1(rst),
    .A2(net48),
    .ZN(_0087_));
 NAND2_X1 _4607_ (.A1(\iir1.y2[9] ),
    .A2(\iir1.y2[10] ),
    .ZN(_0907_));
 XOR2_X1 _4608_ (.A(\iir1.y2[9] ),
    .B(\iir1.y2[7] ),
    .Z(_0908_));
 XNOR2_X1 _4609_ (.A(_0907_),
    .B(_0908_),
    .ZN(_0909_));
 NAND3_X1 _4610_ (.A1(\iir1.y2[8] ),
    .A2(\iir1.y2[6] ),
    .A3(_0909_),
    .ZN(_0910_));
 OAI21_X1 _4611_ (.A(_0910_),
    .B1(_0907_),
    .B2(\iir1.y2[7] ),
    .ZN(_0911_));
 NAND2_X1 _4612_ (.A1(\iir1.y2[8] ),
    .A2(\iir1.y2[6] ),
    .ZN(_0912_));
 XNOR2_X1 _4613_ (.A(_0912_),
    .B(_0909_),
    .ZN(_0913_));
 XOR2_X1 _4614_ (.A(\iir1.y2[9] ),
    .B(\iir1.y2[10] ),
    .Z(_0914_));
 NAND2_X1 _4615_ (.A1(\iir1.y[10] ),
    .A2(_2500_),
    .ZN(_0915_));
 OAI21_X1 _4616_ (.A(_0915_),
    .B1(\iir1.y[10] ),
    .B2(\iir1.y[9] ),
    .ZN(_0916_));
 INV_X1 _4617_ (.A(net45),
    .ZN(_0917_));
 XOR2_X1 _4618_ (.A(\iir1.x1[6] ),
    .B(\iir1.t1[1] ),
    .Z(_0918_));
 NAND3_X1 _4619_ (.A1(\iir1.x1[5] ),
    .A2(\iir1.t1[0] ),
    .A3(_0918_),
    .ZN(_0919_));
 XNOR2_X1 _4620_ (.A(\iir1.x1[7] ),
    .B(\iir1.t1[2] ),
    .ZN(_0920_));
 OR2_X1 _4621_ (.A1(_0919_),
    .A2(_0920_),
    .ZN(_0921_));
 XNOR2_X1 _4622_ (.A(\iir1.x1[8] ),
    .B(\iir1.t1[3] ),
    .ZN(_0922_));
 INV_X1 _4623_ (.A(_0922_),
    .ZN(_0923_));
 NAND2_X1 _4624_ (.A1(\iir1.x1[7] ),
    .A2(\iir1.t1[2] ),
    .ZN(_0924_));
 NAND2_X1 _4625_ (.A1(\iir1.x1[6] ),
    .A2(\iir1.t1[1] ),
    .ZN(_0925_));
 OR2_X1 _4626_ (.A1(_0925_),
    .A2(_0920_),
    .ZN(_0926_));
 NAND2_X1 _4627_ (.A1(_0924_),
    .A2(_0926_),
    .ZN(_0927_));
 XNOR2_X1 _4628_ (.A(_0923_),
    .B(_0927_),
    .ZN(_0928_));
 XNOR2_X1 _4629_ (.A(_0921_),
    .B(_0928_),
    .ZN(_0929_));
 XNOR2_X1 _4630_ (.A(_0917_),
    .B(_0929_),
    .ZN(_0930_));
 XOR2_X1 _4631_ (.A(\iir1.x[5] ),
    .B(_0930_),
    .Z(_0931_));
 NAND2_X1 _4632_ (.A1(_0925_),
    .A2(_0919_),
    .ZN(_0932_));
 XNOR2_X1 _4633_ (.A(_0920_),
    .B(_0932_),
    .ZN(_0933_));
 XNOR2_X1 _4634_ (.A(\iir1.x[5] ),
    .B(_0933_),
    .ZN(_0934_));
 INV_X1 _4635_ (.A(_0934_),
    .ZN(_0935_));
 NAND2_X1 _4636_ (.A1(\iir1.x[4] ),
    .A2(_0935_),
    .ZN(_0936_));
 NAND2_X1 _4637_ (.A1(\iir1.x[5] ),
    .A2(_0933_),
    .ZN(_0937_));
 AOI21_X1 _4638_ (.A(_0931_),
    .B1(_0936_),
    .B2(_0937_),
    .ZN(_0938_));
 AND3_X1 _4639_ (.A1(_0937_),
    .A2(_0936_),
    .A3(_0931_),
    .ZN(_0939_));
 OR2_X1 _4640_ (.A1(_0938_),
    .A2(_0939_),
    .ZN(_0940_));
 INV_X1 _4641_ (.A(_0940_),
    .ZN(_0941_));
 XOR2_X1 _4642_ (.A(\iir1.x[4] ),
    .B(\iir1.x2[6] ),
    .Z(_0942_));
 AOI21_X1 _4643_ (.A(_0938_),
    .B1(_0941_),
    .B2(_0942_),
    .ZN(_0943_));
 NOR2_X1 _4644_ (.A1(_0917_),
    .A2(_0929_),
    .ZN(_0944_));
 INV_X1 _4645_ (.A(_0930_),
    .ZN(_0945_));
 AOI21_X1 _4646_ (.A(_0944_),
    .B1(_0945_),
    .B2(\iir1.x[5] ),
    .ZN(_0946_));
 INV_X1 _4647_ (.A(net43),
    .ZN(_0947_));
 NOR2_X1 _4648_ (.A1(_0921_),
    .A2(_0928_),
    .ZN(_0948_));
 NOR2_X1 _4649_ (.A1(_0926_),
    .A2(_0922_),
    .ZN(_0949_));
 XOR2_X1 _4650_ (.A(\iir1.x1[9] ),
    .B(\iir1.t1[4] ),
    .Z(_0950_));
 NAND2_X1 _4651_ (.A1(\iir1.x1[8] ),
    .A2(\iir1.t1[3] ),
    .ZN(_0951_));
 OAI21_X1 _4652_ (.A(_0951_),
    .B1(_0922_),
    .B2(_0924_),
    .ZN(_0952_));
 XNOR2_X1 _4653_ (.A(_0950_),
    .B(_0952_),
    .ZN(_0953_));
 XNOR2_X1 _4654_ (.A(_0949_),
    .B(_0953_),
    .ZN(_0954_));
 XNOR2_X1 _4655_ (.A(_0948_),
    .B(_0954_),
    .ZN(_0955_));
 XNOR2_X1 _4656_ (.A(_0947_),
    .B(_0955_),
    .ZN(_0956_));
 XNOR2_X1 _4657_ (.A(_0917_),
    .B(_0956_),
    .ZN(_0957_));
 XOR2_X1 _4658_ (.A(_0946_),
    .B(_0957_),
    .Z(_0958_));
 XOR2_X1 _4659_ (.A(\iir1.x[5] ),
    .B(\iir1.x2[7] ),
    .Z(_0959_));
 XNOR2_X1 _4660_ (.A(_0958_),
    .B(_0959_),
    .ZN(_0960_));
 NOR2_X1 _4661_ (.A1(_0943_),
    .A2(_0960_),
    .ZN(_0961_));
 XOR2_X1 _4662_ (.A(_0943_),
    .B(_0960_),
    .Z(_0962_));
 INV_X1 _4663_ (.A(\iir1.x2[6] ),
    .ZN(_0963_));
 OAI211_X1 _4664_ (.A(\iir1.x2[4] ),
    .B(\iir1.x2[5] ),
    .C1(\iir1.x[4] ),
    .C2(_0963_),
    .ZN(_0964_));
 NAND2_X1 _4665_ (.A1(\iir1.x[4] ),
    .A2(\iir1.x2[6] ),
    .ZN(_0965_));
 XNOR2_X1 _4666_ (.A(\iir1.x2[6] ),
    .B(\iir1.x2[5] ),
    .ZN(_0966_));
 XNOR2_X1 _4667_ (.A(_0965_),
    .B(_0966_),
    .ZN(_0967_));
 INV_X1 _4668_ (.A(\iir1.x2[5] ),
    .ZN(_0968_));
 INV_X1 _4669_ (.A(\iir1.x2[4] ),
    .ZN(_0969_));
 OAI21_X1 _4670_ (.A(_0967_),
    .B1(_0968_),
    .B2(_0969_),
    .ZN(_0970_));
 AND2_X1 _4671_ (.A1(_0964_),
    .A2(_0970_),
    .ZN(_0971_));
 AOI21_X1 _4672_ (.A(_0961_),
    .B1(_0962_),
    .B2(_0971_),
    .ZN(_0972_));
 INV_X1 _4673_ (.A(\iir1.x2[7] ),
    .ZN(_0973_));
 OAI211_X1 _4674_ (.A(\iir1.x2[6] ),
    .B(\iir1.x2[5] ),
    .C1(\iir1.x[5] ),
    .C2(_0973_),
    .ZN(_0974_));
 NAND2_X1 _4675_ (.A1(\iir1.x[5] ),
    .A2(\iir1.x2[7] ),
    .ZN(_0975_));
 XNOR2_X1 _4676_ (.A(\iir1.x2[7] ),
    .B(\iir1.x2[6] ),
    .ZN(_0976_));
 XNOR2_X1 _4677_ (.A(_0975_),
    .B(_0976_),
    .ZN(_0977_));
 OAI21_X1 _4678_ (.A(_0977_),
    .B1(_0968_),
    .B2(_0963_),
    .ZN(_0978_));
 AND2_X1 _4679_ (.A1(_0974_),
    .A2(_0978_),
    .ZN(_0979_));
 NOR2_X1 _4680_ (.A1(_0946_),
    .A2(_0957_),
    .ZN(_0980_));
 AOI21_X1 _4681_ (.A(_0980_),
    .B1(_0958_),
    .B2(_0959_),
    .ZN(_0981_));
 XOR2_X1 _4682_ (.A(\iir1.x[6] ),
    .B(\iir1.x2[8] ),
    .Z(_0982_));
 NOR2_X1 _4683_ (.A1(_0947_),
    .A2(_0955_),
    .ZN(_0983_));
 INV_X1 _4684_ (.A(_0956_),
    .ZN(_0984_));
 AOI21_X1 _4685_ (.A(_0983_),
    .B1(_0984_),
    .B2(\iir1.x[6] ),
    .ZN(_0985_));
 NOR3_X1 _4686_ (.A1(_0926_),
    .A2(_0922_),
    .A3(_0953_),
    .ZN(_0986_));
 AOI21_X1 _4687_ (.A(_0986_),
    .B1(_0954_),
    .B2(_0948_),
    .ZN(_0987_));
 NAND4_X1 _4688_ (.A1(\iir1.x1[7] ),
    .A2(\iir1.t1[2] ),
    .A3(_0923_),
    .A4(_0950_),
    .ZN(_0988_));
 XOR2_X1 _4689_ (.A(\iir1.x1[5] ),
    .B(\iir1.x1[10] ),
    .Z(_0989_));
 NAND2_X1 _4690_ (.A1(\iir1.x1[9] ),
    .A2(\iir1.t1[4] ),
    .ZN(_0990_));
 NAND3_X1 _4691_ (.A1(\iir1.x1[8] ),
    .A2(\iir1.t1[3] ),
    .A3(_0950_),
    .ZN(_0991_));
 NAND2_X1 _4692_ (.A1(_0990_),
    .A2(_0991_),
    .ZN(_0992_));
 XOR2_X1 _4693_ (.A(_0989_),
    .B(_0992_),
    .Z(_0993_));
 XOR2_X1 _4694_ (.A(_0988_),
    .B(_0993_),
    .Z(_0994_));
 XOR2_X1 _4695_ (.A(_0987_),
    .B(_0994_),
    .Z(_0995_));
 XNOR2_X1 _4696_ (.A(\iir1.x[8] ),
    .B(_0995_),
    .ZN(_0996_));
 XNOR2_X1 _4697_ (.A(_0947_),
    .B(_0996_),
    .ZN(_0997_));
 XOR2_X1 _4698_ (.A(_0985_),
    .B(_0997_),
    .Z(_0998_));
 XNOR2_X1 _4699_ (.A(_0982_),
    .B(_0998_),
    .ZN(_0999_));
 XOR2_X1 _4700_ (.A(_0981_),
    .B(_0999_),
    .Z(_1000_));
 XNOR2_X1 _4701_ (.A(_0979_),
    .B(_1000_),
    .ZN(_1001_));
 XNOR2_X1 _4702_ (.A(_0972_),
    .B(_1001_),
    .ZN(_1002_));
 OAI21_X1 _4703_ (.A(_0964_),
    .B1(_0965_),
    .B2(\iir1.x2[5] ),
    .ZN(_1003_));
 INV_X1 _4704_ (.A(_1003_),
    .ZN(_1004_));
 OAI22_X1 _4705_ (.A1(_0972_),
    .A2(_1001_),
    .B1(_1002_),
    .B2(_1004_),
    .ZN(_1005_));
 OAI21_X1 _4706_ (.A(_0974_),
    .B1(_0975_),
    .B2(\iir1.x2[6] ),
    .ZN(_1006_));
 NOR2_X1 _4707_ (.A1(_0981_),
    .A2(_0999_),
    .ZN(_1007_));
 AOI21_X1 _4708_ (.A(_1007_),
    .B1(_1000_),
    .B2(_0979_),
    .ZN(_1008_));
 INV_X1 _4709_ (.A(_1008_),
    .ZN(_1009_));
 INV_X1 _4710_ (.A(\iir1.x2[8] ),
    .ZN(_1010_));
 OAI211_X1 _4711_ (.A(\iir1.x2[7] ),
    .B(\iir1.x2[6] ),
    .C1(\iir1.x[6] ),
    .C2(_1010_),
    .ZN(_1011_));
 NAND2_X1 _4712_ (.A1(\iir1.x[6] ),
    .A2(\iir1.x2[8] ),
    .ZN(_1012_));
 XNOR2_X1 _4713_ (.A(\iir1.x2[8] ),
    .B(\iir1.x2[7] ),
    .ZN(_1013_));
 XNOR2_X1 _4714_ (.A(_1012_),
    .B(_1013_),
    .ZN(_1014_));
 OAI21_X1 _4715_ (.A(_1014_),
    .B1(_0963_),
    .B2(_0973_),
    .ZN(_1015_));
 AND2_X1 _4716_ (.A1(_1011_),
    .A2(_1015_),
    .ZN(_1016_));
 NOR2_X1 _4717_ (.A1(_0985_),
    .A2(_0997_),
    .ZN(_1017_));
 AOI21_X1 _4718_ (.A(_1017_),
    .B1(_0998_),
    .B2(_0982_),
    .ZN(_1018_));
 XOR2_X1 _4719_ (.A(\iir1.x[7] ),
    .B(\iir1.x2[9] ),
    .Z(_1019_));
 NOR2_X1 _4720_ (.A1(_0947_),
    .A2(_0996_),
    .ZN(_1020_));
 AOI21_X1 _4721_ (.A(_1020_),
    .B1(_0995_),
    .B2(\iir1.x[8] ),
    .ZN(_1021_));
 INV_X1 _4722_ (.A(net21),
    .ZN(_1022_));
 INV_X1 _4723_ (.A(_0991_),
    .ZN(_1023_));
 NAND2_X1 _4724_ (.A1(_1023_),
    .A2(_0989_),
    .ZN(_1024_));
 NAND3_X1 _4725_ (.A1(\iir1.x1[9] ),
    .A2(\iir1.t1[4] ),
    .A3(_0989_),
    .ZN(_1025_));
 NAND2_X1 _4726_ (.A1(\iir1.x1[5] ),
    .A2(\iir1.x1[10] ),
    .ZN(_1026_));
 XOR2_X1 _4727_ (.A(\iir1.x1[6] ),
    .B(\iir1.x1[10] ),
    .Z(_1027_));
 XNOR2_X1 _4728_ (.A(_1026_),
    .B(_1027_),
    .ZN(_1028_));
 XNOR2_X1 _4729_ (.A(_1025_),
    .B(_1028_),
    .ZN(_1029_));
 XNOR2_X1 _4730_ (.A(_1024_),
    .B(_1029_),
    .ZN(_1030_));
 NOR2_X1 _4731_ (.A1(_0987_),
    .A2(_0994_),
    .ZN(_1031_));
 INV_X1 _4732_ (.A(_0993_),
    .ZN(_1032_));
 NOR2_X1 _4733_ (.A1(_0988_),
    .A2(_1032_),
    .ZN(_1033_));
 OAI21_X1 _4734_ (.A(_1030_),
    .B1(_1031_),
    .B2(_1033_),
    .ZN(_1034_));
 OR3_X1 _4735_ (.A1(_1033_),
    .A2(_1031_),
    .A3(_1030_),
    .ZN(_1035_));
 AND2_X1 _4736_ (.A1(_1034_),
    .A2(_1035_),
    .ZN(_1036_));
 XNOR2_X1 _4737_ (.A(\iir1.x[9] ),
    .B(_1036_),
    .ZN(_1037_));
 XNOR2_X1 _4738_ (.A(_1022_),
    .B(_1037_),
    .ZN(_1038_));
 XOR2_X1 _4739_ (.A(_1021_),
    .B(_1038_),
    .Z(_1039_));
 XNOR2_X1 _4740_ (.A(_1019_),
    .B(_1039_),
    .ZN(_1040_));
 XOR2_X1 _4741_ (.A(_1018_),
    .B(_1040_),
    .Z(_1041_));
 XOR2_X1 _4742_ (.A(_1016_),
    .B(_1041_),
    .Z(_1042_));
 XNOR2_X1 _4743_ (.A(_1009_),
    .B(_1042_),
    .ZN(_1043_));
 XNOR2_X1 _4744_ (.A(_1006_),
    .B(_1043_),
    .ZN(_1044_));
 XNOR2_X1 _4745_ (.A(_1005_),
    .B(_1044_),
    .ZN(_1045_));
 XNOR2_X1 _4746_ (.A(_0962_),
    .B(_0971_),
    .ZN(_1046_));
 XOR2_X1 _4747_ (.A(\iir1.x[4] ),
    .B(_0934_),
    .Z(_1047_));
 NAND2_X1 _4748_ (.A1(\iir1.x1[5] ),
    .A2(\iir1.t1[0] ),
    .ZN(_1048_));
 XNOR2_X1 _4749_ (.A(_1048_),
    .B(_0918_),
    .ZN(_1049_));
 XNOR2_X1 _4750_ (.A(\iir1.x[4] ),
    .B(_1049_),
    .ZN(_1050_));
 INV_X1 _4751_ (.A(_1050_),
    .ZN(_1051_));
 NAND2_X1 _4752_ (.A1(\iir1.x[3] ),
    .A2(_1051_),
    .ZN(_1052_));
 NAND2_X1 _4753_ (.A1(\iir1.x[4] ),
    .A2(_1049_),
    .ZN(_1053_));
 AOI21_X1 _4754_ (.A(_1047_),
    .B1(_1052_),
    .B2(_1053_),
    .ZN(_1054_));
 AND3_X1 _4755_ (.A1(_1053_),
    .A2(_1052_),
    .A3(_1047_),
    .ZN(_1055_));
 OR2_X1 _4756_ (.A1(_1054_),
    .A2(_1055_),
    .ZN(_1056_));
 XNOR2_X1 _4757_ (.A(\iir1.x[3] ),
    .B(\iir1.x2[5] ),
    .ZN(_1057_));
 NOR2_X1 _4758_ (.A1(_1056_),
    .A2(_1057_),
    .ZN(_1058_));
 NOR2_X1 _4759_ (.A1(_1054_),
    .A2(_1058_),
    .ZN(_1059_));
 XNOR2_X1 _4760_ (.A(_0940_),
    .B(_0942_),
    .ZN(_1060_));
 XNOR2_X1 _4761_ (.A(_1059_),
    .B(_1060_),
    .ZN(_1061_));
 NAND2_X1 _4762_ (.A1(\iir1.x2[3] ),
    .A2(\iir1.x2[4] ),
    .ZN(_1062_));
 NAND2_X1 _4763_ (.A1(\iir1.x[3] ),
    .A2(\iir1.x2[5] ),
    .ZN(_1063_));
 XOR2_X1 _4764_ (.A(\iir1.x2[4] ),
    .B(\iir1.x2[5] ),
    .Z(_1064_));
 XNOR2_X1 _4765_ (.A(_1063_),
    .B(_1064_),
    .ZN(_1065_));
 XNOR2_X1 _4766_ (.A(_1062_),
    .B(_1065_),
    .ZN(_1066_));
 NAND2_X1 _4767_ (.A1(_1061_),
    .A2(_1066_),
    .ZN(_1067_));
 OAI21_X1 _4768_ (.A(_1060_),
    .B1(_1058_),
    .B2(_1054_),
    .ZN(_1068_));
 AOI21_X1 _4769_ (.A(_1046_),
    .B1(_1067_),
    .B2(_1068_),
    .ZN(_1069_));
 NAND2_X1 _4770_ (.A1(_1068_),
    .A2(_1067_),
    .ZN(_1070_));
 XNOR2_X1 _4771_ (.A(_1070_),
    .B(_1046_),
    .ZN(_1071_));
 NAND3_X1 _4772_ (.A1(\iir1.x2[3] ),
    .A2(\iir1.x2[4] ),
    .A3(_1065_),
    .ZN(_1072_));
 OAI21_X1 _4773_ (.A(_1072_),
    .B1(_1063_),
    .B2(\iir1.x2[4] ),
    .ZN(_1073_));
 AOI21_X1 _4774_ (.A(_1069_),
    .B1(_1071_),
    .B2(_1073_),
    .ZN(_1074_));
 XNOR2_X1 _4775_ (.A(_1004_),
    .B(_1002_),
    .ZN(_1075_));
 OR2_X1 _4776_ (.A1(_1074_),
    .A2(_1075_),
    .ZN(_1076_));
 XNOR2_X1 _4777_ (.A(_1074_),
    .B(_1075_),
    .ZN(_1077_));
 XNOR2_X1 _4778_ (.A(_1061_),
    .B(_1066_),
    .ZN(_1078_));
 XOR2_X1 _4779_ (.A(\iir1.x[3] ),
    .B(_1050_),
    .Z(_1079_));
 XOR2_X1 _4780_ (.A(\iir1.x1[5] ),
    .B(\iir1.t1[0] ),
    .Z(_1080_));
 XNOR2_X1 _4781_ (.A(\iir1.x[3] ),
    .B(_1080_),
    .ZN(_1081_));
 INV_X1 _4782_ (.A(_1081_),
    .ZN(_1082_));
 NAND2_X1 _4783_ (.A1(\iir1.x[2] ),
    .A2(_1082_),
    .ZN(_1083_));
 NAND2_X1 _4784_ (.A1(\iir1.x[3] ),
    .A2(_1080_),
    .ZN(_1084_));
 AOI21_X1 _4785_ (.A(_1079_),
    .B1(_1083_),
    .B2(_1084_),
    .ZN(_1085_));
 AND3_X1 _4786_ (.A1(_1084_),
    .A2(_1083_),
    .A3(_1079_),
    .ZN(_1086_));
 OR2_X1 _4787_ (.A1(_1085_),
    .A2(_1086_),
    .ZN(_1087_));
 XNOR2_X1 _4788_ (.A(\iir1.x[2] ),
    .B(\iir1.x2[4] ),
    .ZN(_1088_));
 NOR2_X1 _4789_ (.A1(_1087_),
    .A2(_1088_),
    .ZN(_1089_));
 NOR2_X1 _4790_ (.A1(_1085_),
    .A2(_1089_),
    .ZN(_1090_));
 XOR2_X1 _4791_ (.A(_1056_),
    .B(_1057_),
    .Z(_1091_));
 XNOR2_X1 _4792_ (.A(_1090_),
    .B(_1091_),
    .ZN(_1092_));
 NAND2_X1 _4793_ (.A1(\iir1.x2[2] ),
    .A2(\iir1.x2[3] ),
    .ZN(_1093_));
 NAND2_X1 _4794_ (.A1(\iir1.x[2] ),
    .A2(\iir1.x2[4] ),
    .ZN(_1094_));
 XOR2_X1 _4795_ (.A(\iir1.x2[3] ),
    .B(\iir1.x2[4] ),
    .Z(_1095_));
 XNOR2_X1 _4796_ (.A(_1094_),
    .B(_1095_),
    .ZN(_1096_));
 XNOR2_X1 _4797_ (.A(_1093_),
    .B(_1096_),
    .ZN(_1097_));
 NAND2_X1 _4798_ (.A1(_1092_),
    .A2(_1097_),
    .ZN(_1098_));
 OAI21_X1 _4799_ (.A(_1091_),
    .B1(_1089_),
    .B2(_1085_),
    .ZN(_1099_));
 AOI21_X1 _4800_ (.A(_1078_),
    .B1(_1098_),
    .B2(_1099_),
    .ZN(_1100_));
 NAND2_X1 _4801_ (.A1(_1099_),
    .A2(_1098_),
    .ZN(_1101_));
 XNOR2_X1 _4802_ (.A(_1101_),
    .B(_1078_),
    .ZN(_1102_));
 NAND3_X1 _4803_ (.A1(\iir1.x2[2] ),
    .A2(\iir1.x2[3] ),
    .A3(_1096_),
    .ZN(_1103_));
 OAI21_X1 _4804_ (.A(_1103_),
    .B1(_1094_),
    .B2(\iir1.x2[3] ),
    .ZN(_1104_));
 AOI21_X1 _4805_ (.A(_1100_),
    .B1(_1102_),
    .B2(_1104_),
    .ZN(_1105_));
 XNOR2_X1 _4806_ (.A(_1071_),
    .B(_1073_),
    .ZN(_1106_));
 NOR2_X1 _4807_ (.A1(_1105_),
    .A2(_1106_),
    .ZN(_1107_));
 XOR2_X1 _4808_ (.A(_1105_),
    .B(_1106_),
    .Z(_1108_));
 AND2_X1 _4809_ (.A1(\iir1.t1[4] ),
    .A2(\iir1.x[2] ),
    .ZN(_1109_));
 XOR2_X1 _4810_ (.A(\iir1.t1[4] ),
    .B(\iir1.x[2] ),
    .Z(_1110_));
 AOI21_X1 _4811_ (.A(_1109_),
    .B1(_1110_),
    .B2(\iir1.x[1] ),
    .ZN(_1111_));
 XOR2_X1 _4812_ (.A(\iir1.x[2] ),
    .B(_1081_),
    .Z(_1112_));
 XOR2_X1 _4813_ (.A(_1111_),
    .B(_1112_),
    .Z(_1113_));
 XOR2_X1 _4814_ (.A(\iir1.x[1] ),
    .B(\iir1.x2[3] ),
    .Z(_1114_));
 NAND2_X1 _4815_ (.A1(_1113_),
    .A2(_1114_),
    .ZN(_1115_));
 OAI21_X1 _4816_ (.A(_1115_),
    .B1(_1112_),
    .B2(_1111_),
    .ZN(_1116_));
 XOR2_X1 _4817_ (.A(_1087_),
    .B(_1088_),
    .Z(_1117_));
 XOR2_X1 _4818_ (.A(_1116_),
    .B(_1117_),
    .Z(_1118_));
 NAND2_X1 _4819_ (.A1(\iir1.x2[1] ),
    .A2(\iir1.x2[2] ),
    .ZN(_1119_));
 NAND2_X1 _4820_ (.A1(\iir1.x[1] ),
    .A2(\iir1.x2[3] ),
    .ZN(_1120_));
 XOR2_X1 _4821_ (.A(\iir1.x2[2] ),
    .B(\iir1.x2[3] ),
    .Z(_1121_));
 XNOR2_X1 _4822_ (.A(_1120_),
    .B(_1121_),
    .ZN(_1122_));
 XNOR2_X1 _4823_ (.A(_1119_),
    .B(_1122_),
    .ZN(_1123_));
 AOI22_X1 _4824_ (.A1(_1116_),
    .A2(_1117_),
    .B1(_1118_),
    .B2(_1123_),
    .ZN(_1124_));
 XNOR2_X1 _4825_ (.A(_1092_),
    .B(_1097_),
    .ZN(_1125_));
 XOR2_X1 _4826_ (.A(_1124_),
    .B(_1125_),
    .Z(_1126_));
 NAND3_X1 _4827_ (.A1(\iir1.x2[1] ),
    .A2(\iir1.x2[2] ),
    .A3(_1122_),
    .ZN(_1127_));
 OAI21_X1 _4828_ (.A(_1127_),
    .B1(_1120_),
    .B2(\iir1.x2[2] ),
    .ZN(_1128_));
 NAND2_X1 _4829_ (.A1(_1126_),
    .A2(_1128_),
    .ZN(_1129_));
 OAI21_X1 _4830_ (.A(_1129_),
    .B1(_1125_),
    .B2(_1124_),
    .ZN(_1130_));
 XOR2_X1 _4831_ (.A(_1102_),
    .B(_1104_),
    .Z(_1131_));
 NAND2_X1 _4832_ (.A1(_1130_),
    .A2(_1131_),
    .ZN(_1132_));
 XNOR2_X1 _4833_ (.A(_1126_),
    .B(_1128_),
    .ZN(_1133_));
 XNOR2_X1 _4834_ (.A(\iir1.x[1] ),
    .B(_1110_),
    .ZN(_1134_));
 NOR2_X1 _4835_ (.A1(\iir1.t1[3] ),
    .A2(\iir1.x[1] ),
    .ZN(_1135_));
 AOI21_X1 _4836_ (.A(\iir1.x[0] ),
    .B1(\iir1.x[1] ),
    .B2(\iir1.t1[3] ),
    .ZN(_1136_));
 NOR3_X1 _4837_ (.A1(_1134_),
    .A2(_1135_),
    .A3(_1136_),
    .ZN(_1137_));
 NOR2_X1 _4838_ (.A1(_1135_),
    .A2(_1136_),
    .ZN(_1138_));
 XNOR2_X1 _4839_ (.A(_1134_),
    .B(_1138_),
    .ZN(_1139_));
 XOR2_X1 _4840_ (.A(\iir1.x[0] ),
    .B(\iir1.x2[2] ),
    .Z(_1140_));
 AOI21_X1 _4841_ (.A(_1137_),
    .B1(_1139_),
    .B2(_1140_),
    .ZN(_1141_));
 XNOR2_X1 _4842_ (.A(_1113_),
    .B(_1114_),
    .ZN(_1142_));
 NOR2_X1 _4843_ (.A1(_1141_),
    .A2(_1142_),
    .ZN(_1143_));
 XOR2_X1 _4844_ (.A(_1141_),
    .B(_1142_),
    .Z(_1144_));
 NAND2_X1 _4845_ (.A1(\iir1.x2[0] ),
    .A2(\iir1.x2[1] ),
    .ZN(_1145_));
 NAND2_X1 _4846_ (.A1(\iir1.x[0] ),
    .A2(\iir1.x2[2] ),
    .ZN(_1146_));
 XOR2_X1 _4847_ (.A(\iir1.x2[1] ),
    .B(\iir1.x2[2] ),
    .Z(_1147_));
 XNOR2_X1 _4848_ (.A(_1146_),
    .B(_1147_),
    .ZN(_1148_));
 XNOR2_X1 _4849_ (.A(_1145_),
    .B(_1148_),
    .ZN(_1149_));
 AOI21_X1 _4850_ (.A(_1143_),
    .B1(_1144_),
    .B2(_1149_),
    .ZN(_1150_));
 XNOR2_X1 _4851_ (.A(_1118_),
    .B(_1123_),
    .ZN(_1151_));
 XOR2_X1 _4852_ (.A(_1150_),
    .B(_1151_),
    .Z(_1152_));
 AOI21_X1 _4853_ (.A(_1147_),
    .B1(\iir1.x2[2] ),
    .B2(\iir1.x[0] ),
    .ZN(_1153_));
 OAI22_X1 _4854_ (.A1(\iir1.x2[1] ),
    .A2(_1146_),
    .B1(_1145_),
    .B2(_1153_),
    .ZN(_1154_));
 NAND2_X1 _4855_ (.A1(_1152_),
    .A2(_1154_),
    .ZN(_1155_));
 OR2_X1 _4856_ (.A1(_1150_),
    .A2(_1151_),
    .ZN(_1156_));
 AOI21_X1 _4857_ (.A(_1133_),
    .B1(_1155_),
    .B2(_1156_),
    .ZN(_1157_));
 NAND2_X1 _4858_ (.A1(_1156_),
    .A2(_1155_),
    .ZN(_1158_));
 XNOR2_X1 _4859_ (.A(_1158_),
    .B(_1133_),
    .ZN(_1159_));
 XNOR2_X1 _4860_ (.A(_1144_),
    .B(_1149_),
    .ZN(_1160_));
 XOR2_X1 _4861_ (.A(\iir1.t1[3] ),
    .B(\iir1.x[1] ),
    .Z(_1161_));
 INV_X1 _4862_ (.A(net6),
    .ZN(_1162_));
 NAND2_X1 _4863_ (.A1(_1162_),
    .A2(\iir1.x[0] ),
    .ZN(_1163_));
 XNOR2_X1 _4864_ (.A(_1161_),
    .B(_1163_),
    .ZN(_1164_));
 NAND2_X1 _4865_ (.A1(\iir1.x2[1] ),
    .A2(_1164_),
    .ZN(_1165_));
 NAND2_X1 _4866_ (.A1(\iir1.t1[2] ),
    .A2(\iir1.x[0] ),
    .ZN(_1166_));
 OAI21_X1 _4867_ (.A(_1165_),
    .B1(_1166_),
    .B2(_1161_),
    .ZN(_1167_));
 XNOR2_X1 _4868_ (.A(_1139_),
    .B(_1140_),
    .ZN(_1168_));
 INV_X1 _4869_ (.A(_1168_),
    .ZN(_1169_));
 XNOR2_X1 _4870_ (.A(_1167_),
    .B(_1169_),
    .ZN(_1170_));
 XNOR2_X1 _4871_ (.A(\iir1.x2[0] ),
    .B(\iir1.x2[1] ),
    .ZN(_1171_));
 OR2_X1 _4872_ (.A1(_1170_),
    .A2(_1171_),
    .ZN(_1172_));
 NAND2_X1 _4873_ (.A1(_1167_),
    .A2(_1169_),
    .ZN(_1173_));
 AOI21_X1 _4874_ (.A(_1160_),
    .B1(_1172_),
    .B2(_1173_),
    .ZN(_1174_));
 XOR2_X1 _4875_ (.A(_1152_),
    .B(_1154_),
    .Z(_1175_));
 NAND2_X1 _4876_ (.A1(_1174_),
    .A2(_1175_),
    .ZN(_1176_));
 INV_X1 _4877_ (.A(\iir1.x2[0] ),
    .ZN(_1177_));
 XOR2_X1 _4878_ (.A(\iir1.t1[2] ),
    .B(\iir1.x[0] ),
    .Z(_1178_));
 NAND2_X1 _4879_ (.A1(\iir1.x2[0] ),
    .A2(_1178_),
    .ZN(_1179_));
 XNOR2_X1 _4880_ (.A(\iir1.x2[1] ),
    .B(_1164_),
    .ZN(_1180_));
 AOI21_X1 _4881_ (.A(_1177_),
    .B1(_1179_),
    .B2(_1180_),
    .ZN(_1181_));
 XOR2_X1 _4882_ (.A(_1170_),
    .B(_1171_),
    .Z(_1182_));
 AND3_X1 _4883_ (.A1(_1173_),
    .A2(_1172_),
    .A3(_1160_),
    .ZN(_1183_));
 NOR2_X1 _4884_ (.A1(_1174_),
    .A2(_1183_),
    .ZN(_1184_));
 NAND3_X1 _4885_ (.A1(_1181_),
    .A2(_1182_),
    .A3(_1184_),
    .ZN(_1185_));
 XNOR2_X1 _4886_ (.A(_1174_),
    .B(_1175_),
    .ZN(_1186_));
 OAI21_X1 _4887_ (.A(_1176_),
    .B1(_1185_),
    .B2(_1186_),
    .ZN(_1187_));
 AOI21_X1 _4888_ (.A(_1157_),
    .B1(_1159_),
    .B2(_1187_),
    .ZN(_1188_));
 NOR2_X1 _4889_ (.A1(_1130_),
    .A2(_1131_),
    .ZN(_1189_));
 OAI21_X1 _4890_ (.A(_1132_),
    .B1(_1188_),
    .B2(_1189_),
    .ZN(_1190_));
 AOI21_X1 _4891_ (.A(_1107_),
    .B1(_1108_),
    .B2(_1190_),
    .ZN(_1191_));
 OAI21_X1 _4892_ (.A(_1076_),
    .B1(_1077_),
    .B2(_1191_),
    .ZN(_1192_));
 XOR2_X1 _4893_ (.A(_1045_),
    .B(_1192_),
    .Z(_1193_));
 XNOR2_X1 _4894_ (.A(\iir1.y[1] ),
    .B(_1193_),
    .ZN(_1194_));
 XNOR2_X1 _4895_ (.A(_1191_),
    .B(_1077_),
    .ZN(_1195_));
 NOR2_X1 _4896_ (.A1(_0006_),
    .A2(_1195_),
    .ZN(_1196_));
 XOR2_X1 _4897_ (.A(\iir1.y[10] ),
    .B(_1195_),
    .Z(_1197_));
 NOR2_X1 _4898_ (.A1(_0737_),
    .A2(_1197_),
    .ZN(_1198_));
 OAI21_X1 _4899_ (.A(_1194_),
    .B1(_1196_),
    .B2(_1198_),
    .ZN(_1199_));
 OR3_X1 _4900_ (.A1(_1198_),
    .A2(_1196_),
    .A3(_1194_),
    .ZN(_1200_));
 AND2_X1 _4901_ (.A1(_1199_),
    .A2(_1200_),
    .ZN(_1201_));
 NAND2_X1 _4902_ (.A1(\iir1.y[2] ),
    .A2(_1201_),
    .ZN(_1202_));
 NAND2_X1 _4903_ (.A1(_1199_),
    .A2(_1202_),
    .ZN(_1203_));
 NAND2_X1 _4904_ (.A1(_1572_),
    .A2(_1627_),
    .ZN(_1204_));
 INV_X1 _4905_ (.A(_1193_),
    .ZN(_1205_));
 NAND2_X1 _4906_ (.A1(\iir1.y[1] ),
    .A2(_1205_),
    .ZN(_1206_));
 NAND2_X1 _4907_ (.A1(_1005_),
    .A2(_1044_),
    .ZN(_1207_));
 OR3_X1 _4908_ (.A1(_1191_),
    .A2(_1077_),
    .A3(_1045_),
    .ZN(_1208_));
 OAI211_X1 _4909_ (.A(_1207_),
    .B(_1208_),
    .C1(_1045_),
    .C2(_1076_),
    .ZN(_1209_));
 INV_X1 _4910_ (.A(_1043_),
    .ZN(_1210_));
 AOI22_X1 _4911_ (.A1(_1009_),
    .A2(_1042_),
    .B1(_1210_),
    .B2(_1006_),
    .ZN(_1211_));
 OAI21_X1 _4912_ (.A(_1011_),
    .B1(_1012_),
    .B2(\iir1.x2[7] ),
    .ZN(_1212_));
 INV_X1 _4913_ (.A(_1212_),
    .ZN(_1213_));
 NOR2_X1 _4914_ (.A1(_1018_),
    .A2(_1040_),
    .ZN(_1214_));
 AOI21_X1 _4915_ (.A(_1214_),
    .B1(_1041_),
    .B2(_1016_),
    .ZN(_1215_));
 INV_X1 _4916_ (.A(\iir1.x2[9] ),
    .ZN(_1216_));
 OAI211_X1 _4917_ (.A(\iir1.x2[8] ),
    .B(\iir1.x2[7] ),
    .C1(\iir1.x[7] ),
    .C2(_1216_),
    .ZN(_1217_));
 NAND2_X1 _4918_ (.A1(\iir1.x[7] ),
    .A2(\iir1.x2[9] ),
    .ZN(_1218_));
 XNOR2_X1 _4919_ (.A(\iir1.x2[9] ),
    .B(\iir1.x2[8] ),
    .ZN(_1219_));
 XNOR2_X1 _4920_ (.A(_1218_),
    .B(_1219_),
    .ZN(_1220_));
 OAI21_X1 _4921_ (.A(_1220_),
    .B1(_0973_),
    .B2(_1010_),
    .ZN(_1221_));
 AND2_X1 _4922_ (.A1(_1217_),
    .A2(_1221_),
    .ZN(_1222_));
 NOR2_X1 _4923_ (.A1(_1021_),
    .A2(_1038_),
    .ZN(_1223_));
 AOI21_X1 _4924_ (.A(_1223_),
    .B1(_1039_),
    .B2(_1019_),
    .ZN(_1224_));
 XOR2_X1 _4925_ (.A(\iir1.x[8] ),
    .B(\iir1.x2[10] ),
    .Z(_1225_));
 INV_X1 _4926_ (.A(_1225_),
    .ZN(_1226_));
 NAND2_X1 _4927_ (.A1(\iir1.x[9] ),
    .A2(_1036_),
    .ZN(_1227_));
 OAI21_X1 _4928_ (.A(_1227_),
    .B1(_1037_),
    .B2(_1022_),
    .ZN(_1228_));
 INV_X1 _4929_ (.A(_1228_),
    .ZN(_1229_));
 INV_X1 _4930_ (.A(net24),
    .ZN(_1230_));
 NAND3_X1 _4931_ (.A1(_1023_),
    .A2(_0989_),
    .A3(_1029_),
    .ZN(_1231_));
 AND4_X1 _4932_ (.A1(\iir1.x1[9] ),
    .A2(\iir1.t1[4] ),
    .A3(_0989_),
    .A4(_1028_),
    .ZN(_1232_));
 INV_X1 _4933_ (.A(net1),
    .ZN(_1233_));
 NAND2_X1 _4934_ (.A1(_1233_),
    .A2(\iir1.x1[10] ),
    .ZN(_1234_));
 OR3_X1 _4935_ (.A1(\iir1.x1[7] ),
    .A2(\iir1.x1[5] ),
    .A3(_1234_),
    .ZN(_1235_));
 OAI21_X1 _4936_ (.A(\iir1.x1[7] ),
    .B1(\iir1.x1[5] ),
    .B2(_1234_),
    .ZN(_1236_));
 AND2_X1 _4937_ (.A1(_1235_),
    .A2(_1236_),
    .ZN(_1237_));
 XOR2_X1 _4938_ (.A(_1232_),
    .B(_1237_),
    .Z(_1238_));
 AND3_X1 _4939_ (.A1(_1231_),
    .A2(_1034_),
    .A3(_1238_),
    .ZN(_1239_));
 AOI21_X1 _4940_ (.A(_1238_),
    .B1(_1034_),
    .B2(_1231_),
    .ZN(_1240_));
 OR2_X1 _4941_ (.A1(_1239_),
    .A2(_1240_),
    .ZN(_1241_));
 XOR2_X1 _4942_ (.A(\iir1.x[10] ),
    .B(_1241_),
    .Z(_1242_));
 XNOR2_X1 _4943_ (.A(_1230_),
    .B(_1242_),
    .ZN(_1243_));
 XNOR2_X1 _4944_ (.A(_1229_),
    .B(_1243_),
    .ZN(_1244_));
 XNOR2_X1 _4945_ (.A(_1226_),
    .B(_1244_),
    .ZN(_1245_));
 XOR2_X1 _4946_ (.A(_1224_),
    .B(_1245_),
    .Z(_1246_));
 XNOR2_X1 _4947_ (.A(_1222_),
    .B(_1246_),
    .ZN(_1247_));
 XNOR2_X1 _4948_ (.A(_1215_),
    .B(_1247_),
    .ZN(_1248_));
 XNOR2_X1 _4949_ (.A(_1213_),
    .B(_1248_),
    .ZN(_1249_));
 XOR2_X1 _4950_ (.A(_1211_),
    .B(_1249_),
    .Z(_1250_));
 XNOR2_X1 _4951_ (.A(_1209_),
    .B(_1250_),
    .ZN(_1251_));
 XOR2_X1 _4952_ (.A(_1206_),
    .B(_1251_),
    .Z(_1252_));
 XNOR2_X1 _4953_ (.A(_1204_),
    .B(_1252_),
    .ZN(_1253_));
 XNOR2_X1 _4954_ (.A(_1203_),
    .B(_1253_),
    .ZN(_1254_));
 XNOR2_X1 _4955_ (.A(\iir1.y[7] ),
    .B(_1254_),
    .ZN(_1255_));
 XNOR2_X1 _4956_ (.A(\iir1.y[2] ),
    .B(_1201_),
    .ZN(_1256_));
 XNOR2_X1 _4957_ (.A(_1190_),
    .B(_1108_),
    .ZN(_1257_));
 NAND2_X1 _4958_ (.A1(\iir1.y[0] ),
    .A2(_1257_),
    .ZN(_1258_));
 XOR2_X1 _4959_ (.A(_1197_),
    .B(_1258_),
    .Z(_1259_));
 NAND2_X1 _4960_ (.A1(\iir1.y[1] ),
    .A2(_1259_),
    .ZN(_1260_));
 INV_X1 _4961_ (.A(_1257_),
    .ZN(_1261_));
 NAND3_X1 _4962_ (.A1(\iir1.y[0] ),
    .A2(_1261_),
    .A3(_1197_),
    .ZN(_1262_));
 AOI21_X1 _4963_ (.A(_1256_),
    .B1(_1260_),
    .B2(_1262_),
    .ZN(_1263_));
 AND3_X1 _4964_ (.A1(_1262_),
    .A2(_1260_),
    .A3(_1256_),
    .ZN(_1264_));
 NOR2_X1 _4965_ (.A1(_1263_),
    .A2(_1264_),
    .ZN(_1265_));
 AND2_X1 _4966_ (.A1(\iir1.y[6] ),
    .A2(_1265_),
    .ZN(_1266_));
 OAI21_X1 _4967_ (.A(_1255_),
    .B1(_1266_),
    .B2(_1263_),
    .ZN(_1267_));
 OR3_X1 _4968_ (.A1(_1263_),
    .A2(_1266_),
    .A3(_1255_),
    .ZN(_1268_));
 AND2_X1 _4969_ (.A1(_1267_),
    .A2(_1268_),
    .ZN(_1269_));
 XOR2_X1 _4970_ (.A(_0916_),
    .B(_1269_),
    .Z(_1270_));
 NOR2_X1 _4971_ (.A1(\iir1.y[8] ),
    .A2(\iir1.y[10] ),
    .ZN(_1271_));
 NOR2_X1 _4972_ (.A1(_2647_),
    .A2(_1271_),
    .ZN(_1272_));
 XNOR2_X1 _4973_ (.A(_0737_),
    .B(_1257_),
    .ZN(_1273_));
 INV_X1 _4974_ (.A(_1273_),
    .ZN(_1274_));
 NAND2_X1 _4975_ (.A1(\iir1.y[4] ),
    .A2(_1274_),
    .ZN(_1275_));
 XNOR2_X1 _4976_ (.A(\iir1.y[1] ),
    .B(_1259_),
    .ZN(_1276_));
 NOR2_X1 _4977_ (.A1(_1275_),
    .A2(_1276_),
    .ZN(_1277_));
 XOR2_X1 _4978_ (.A(_1275_),
    .B(_1276_),
    .Z(_1278_));
 AOI21_X1 _4979_ (.A(_1277_),
    .B1(_1278_),
    .B2(\iir1.y[5] ),
    .ZN(_1279_));
 XNOR2_X1 _4980_ (.A(\iir1.y[6] ),
    .B(_1265_),
    .ZN(_1280_));
 XOR2_X1 _4981_ (.A(_1279_),
    .B(_1280_),
    .Z(_1281_));
 NAND2_X1 _4982_ (.A1(_1272_),
    .A2(_1281_),
    .ZN(_1282_));
 OR2_X1 _4983_ (.A1(_1279_),
    .A2(_1280_),
    .ZN(_1283_));
 AOI21_X1 _4984_ (.A(_1270_),
    .B1(_1282_),
    .B2(_1283_),
    .ZN(_1284_));
 NAND2_X1 _4985_ (.A1(_1203_),
    .A2(_1253_),
    .ZN(_1285_));
 INV_X1 _4986_ (.A(net94),
    .ZN(_1286_));
 OAI21_X1 _4987_ (.A(_1285_),
    .B1(_1254_),
    .B2(_1286_),
    .ZN(_1287_));
 NAND3_X1 _4988_ (.A1(_1572_),
    .A2(_1627_),
    .A3(_1252_),
    .ZN(_1288_));
 OAI21_X1 _4989_ (.A(_1288_),
    .B1(_1251_),
    .B2(_1206_),
    .ZN(_1289_));
 NOR2_X1 _4990_ (.A1(_1211_),
    .A2(_1249_),
    .ZN(_1290_));
 AOI21_X1 _4991_ (.A(_1290_),
    .B1(_1250_),
    .B2(_1209_),
    .ZN(_1291_));
 OAI21_X1 _4992_ (.A(_1217_),
    .B1(_1218_),
    .B2(\iir1.x2[8] ),
    .ZN(_1292_));
 NOR2_X1 _4993_ (.A1(_1224_),
    .A2(_1245_),
    .ZN(_1293_));
 AOI21_X1 _4994_ (.A(_1293_),
    .B1(_1246_),
    .B2(_1222_),
    .ZN(_1294_));
 INV_X1 _4995_ (.A(\iir1.x2[10] ),
    .ZN(_1295_));
 OAI211_X1 _4996_ (.A(\iir1.x2[9] ),
    .B(\iir1.x2[8] ),
    .C1(\iir1.x[8] ),
    .C2(_1295_),
    .ZN(_1296_));
 NAND2_X1 _4997_ (.A1(\iir1.x[8] ),
    .A2(\iir1.x2[10] ),
    .ZN(_1298_));
 XNOR2_X1 _4998_ (.A(\iir1.x2[10] ),
    .B(\iir1.x2[9] ),
    .ZN(_1299_));
 XNOR2_X1 _4999_ (.A(_1298_),
    .B(_1299_),
    .ZN(_1300_));
 OAI21_X1 _5000_ (.A(_1300_),
    .B1(_1010_),
    .B2(_1216_),
    .ZN(_1301_));
 AND2_X1 _5001_ (.A1(_1296_),
    .A2(_1301_),
    .ZN(_1302_));
 OR2_X1 _5002_ (.A1(_1229_),
    .A2(_1243_),
    .ZN(_1303_));
 OAI21_X1 _5003_ (.A(_1303_),
    .B1(_1244_),
    .B2(_1226_),
    .ZN(_1304_));
 XNOR2_X1 _5004_ (.A(\iir1.x[9] ),
    .B(\iir1.x2[10] ),
    .ZN(_1305_));
 OAI22_X1 _5005_ (.A1(_0010_),
    .A2(_1241_),
    .B1(_1242_),
    .B2(_1230_),
    .ZN(_1306_));
 NOR3_X1 _5006_ (.A1(\iir1.x1[8] ),
    .A2(\iir1.x1[7] ),
    .A3(_1234_),
    .ZN(_1307_));
 AOI21_X1 _5007_ (.A(_1307_),
    .B1(_1235_),
    .B2(\iir1.x1[8] ),
    .ZN(_1309_));
 AOI21_X1 _5008_ (.A(_1309_),
    .B1(_1307_),
    .B2(\iir1.x1[5] ),
    .ZN(_1310_));
 INV_X1 _5009_ (.A(_1237_),
    .ZN(_1311_));
 AOI21_X1 _5010_ (.A(_1240_),
    .B1(_1311_),
    .B2(_1232_),
    .ZN(_1312_));
 XNOR2_X1 _5011_ (.A(_1310_),
    .B(_1312_),
    .ZN(_1313_));
 XNOR2_X1 _5012_ (.A(_1306_),
    .B(_1313_),
    .ZN(_1314_));
 XOR2_X1 _5013_ (.A(_1305_),
    .B(_1314_),
    .Z(_1315_));
 XOR2_X1 _5014_ (.A(_1304_),
    .B(_1315_),
    .Z(_1316_));
 XNOR2_X1 _5015_ (.A(_1302_),
    .B(_1316_),
    .ZN(_1317_));
 XNOR2_X1 _5016_ (.A(_1294_),
    .B(_1317_),
    .ZN(_1318_));
 XNOR2_X1 _5017_ (.A(_1292_),
    .B(_1318_),
    .ZN(_1320_));
 NOR2_X1 _5018_ (.A1(_1213_),
    .A2(_1248_),
    .ZN(_1321_));
 OR2_X1 _5019_ (.A1(_1215_),
    .A2(_1247_),
    .ZN(_1322_));
 INV_X1 _5020_ (.A(_1322_),
    .ZN(_1323_));
 OAI21_X1 _5021_ (.A(_1320_),
    .B1(_1321_),
    .B2(_1323_),
    .ZN(_1324_));
 OR3_X1 _5022_ (.A1(_1323_),
    .A2(_1321_),
    .A3(_1320_),
    .ZN(_1325_));
 NAND2_X1 _5023_ (.A1(_1324_),
    .A2(_1325_),
    .ZN(_1326_));
 XOR2_X1 _5024_ (.A(_1291_),
    .B(_1326_),
    .Z(_1327_));
 XOR2_X1 _5025_ (.A(_1550_),
    .B(_1327_),
    .Z(_1328_));
 XNOR2_X1 _5026_ (.A(_1289_),
    .B(_1328_),
    .ZN(_1329_));
 XOR2_X1 _5027_ (.A(_1572_),
    .B(_1329_),
    .Z(_1331_));
 XNOR2_X1 _5028_ (.A(_1287_),
    .B(_1331_),
    .ZN(_1332_));
 XOR2_X1 _5029_ (.A(_0005_),
    .B(_2722_),
    .Z(_1333_));
 XNOR2_X1 _5030_ (.A(_1332_),
    .B(_1333_),
    .ZN(_1334_));
 OAI211_X1 _5031_ (.A(_0915_),
    .B(_1269_),
    .C1(\iir1.y[9] ),
    .C2(\iir1.y[10] ),
    .ZN(_1335_));
 AOI21_X1 _5032_ (.A(_1334_),
    .B1(_1335_),
    .B2(_1267_),
    .ZN(_1336_));
 AND3_X1 _5033_ (.A1(_1267_),
    .A2(_1335_),
    .A3(_1334_),
    .ZN(_1337_));
 NOR2_X1 _5034_ (.A1(_1336_),
    .A2(_1337_),
    .ZN(_1338_));
 AND2_X1 _5035_ (.A1(_1284_),
    .A2(_1338_),
    .ZN(_1339_));
 XOR2_X1 _5036_ (.A(_1284_),
    .B(_1338_),
    .Z(_1340_));
 XNOR2_X1 _5037_ (.A(_1272_),
    .B(_1281_),
    .ZN(_1342_));
 XOR2_X1 _5038_ (.A(_1130_),
    .B(_1131_),
    .Z(_1343_));
 XNOR2_X1 _5039_ (.A(_1188_),
    .B(_1343_),
    .ZN(_1344_));
 NAND2_X1 _5040_ (.A1(\iir1.y[3] ),
    .A2(_1344_),
    .ZN(_1345_));
 XOR2_X1 _5041_ (.A(\iir1.y[4] ),
    .B(_1273_),
    .Z(_1346_));
 NOR2_X1 _5042_ (.A1(_1345_),
    .A2(_1346_),
    .ZN(_1347_));
 XOR2_X1 _5043_ (.A(_1345_),
    .B(_1346_),
    .Z(_1348_));
 AOI21_X1 _5044_ (.A(_1347_),
    .B1(_1348_),
    .B2(\iir1.y[6] ),
    .ZN(_1349_));
 XNOR2_X1 _5045_ (.A(\iir1.y[5] ),
    .B(_1278_),
    .ZN(_1350_));
 XOR2_X1 _5046_ (.A(_1349_),
    .B(_1350_),
    .Z(_1351_));
 NAND2_X1 _5047_ (.A1(\iir1.y[7] ),
    .A2(_1351_),
    .ZN(_1353_));
 OR2_X1 _5048_ (.A1(_1349_),
    .A2(_1350_),
    .ZN(_1354_));
 AOI21_X1 _5049_ (.A(_1342_),
    .B1(_1353_),
    .B2(_1354_),
    .ZN(_1355_));
 AND3_X1 _5050_ (.A1(_1283_),
    .A2(_1282_),
    .A3(_1270_),
    .ZN(_1356_));
 NOR2_X1 _5051_ (.A1(_1284_),
    .A2(_1356_),
    .ZN(_1357_));
 NAND2_X1 _5052_ (.A1(_1355_),
    .A2(_1357_),
    .ZN(_1358_));
 XNOR2_X1 _5053_ (.A(_1355_),
    .B(_1357_),
    .ZN(_1359_));
 NAND2_X1 _5054_ (.A1(_1354_),
    .A2(_1353_),
    .ZN(_1360_));
 XNOR2_X1 _5055_ (.A(_1360_),
    .B(_1342_),
    .ZN(_1361_));
 NOR3_X1 _5056_ (.A1(_0000_),
    .A2(_0007_),
    .A3(_2436_),
    .ZN(_1362_));
 XNOR2_X1 _5057_ (.A(\iir1.y[7] ),
    .B(_1351_),
    .ZN(_1364_));
 XOR2_X1 _5058_ (.A(_1185_),
    .B(_1186_),
    .Z(_1365_));
 AND2_X1 _5059_ (.A1(\iir1.y[1] ),
    .A2(_1365_),
    .ZN(_1366_));
 XOR2_X1 _5060_ (.A(_1159_),
    .B(_1187_),
    .Z(_1367_));
 NAND2_X1 _5061_ (.A1(_1366_),
    .A2(_1367_),
    .ZN(_1368_));
 NOR2_X1 _5062_ (.A1(_1366_),
    .A2(_1367_),
    .ZN(_1369_));
 OAI21_X1 _5063_ (.A(_1368_),
    .B1(_1369_),
    .B2(_2336_),
    .ZN(_1370_));
 INV_X1 _5064_ (.A(_1370_),
    .ZN(_1371_));
 XNOR2_X1 _5065_ (.A(\iir1.y[3] ),
    .B(_1344_),
    .ZN(_1372_));
 NOR2_X1 _5066_ (.A1(_1371_),
    .A2(_1372_),
    .ZN(_1373_));
 NAND2_X1 _5067_ (.A1(_1371_),
    .A2(_1372_),
    .ZN(_1375_));
 XOR2_X1 _5068_ (.A(_0007_),
    .B(_2436_),
    .Z(_1376_));
 AOI21_X1 _5069_ (.A(_1373_),
    .B1(_1375_),
    .B2(_1376_),
    .ZN(_1377_));
 XNOR2_X1 _5070_ (.A(\iir1.y[6] ),
    .B(_1348_),
    .ZN(_1378_));
 XOR2_X1 _5071_ (.A(_1377_),
    .B(_1378_),
    .Z(_1379_));
 NOR2_X1 _5072_ (.A1(_0007_),
    .A2(_2436_),
    .ZN(_1380_));
 XNOR2_X1 _5073_ (.A(_0000_),
    .B(_1380_),
    .ZN(_1381_));
 NAND2_X1 _5074_ (.A1(_1379_),
    .A2(_1381_),
    .ZN(_1382_));
 OR2_X1 _5075_ (.A1(_1377_),
    .A2(_1378_),
    .ZN(_1383_));
 AOI21_X1 _5076_ (.A(_1364_),
    .B1(_1382_),
    .B2(_1383_),
    .ZN(_1384_));
 AND3_X1 _5077_ (.A1(_1383_),
    .A2(_1382_),
    .A3(_1364_),
    .ZN(_1386_));
 NOR2_X1 _5078_ (.A1(_1384_),
    .A2(_1386_),
    .ZN(_1387_));
 AND2_X1 _5079_ (.A1(_1362_),
    .A2(_1387_),
    .ZN(_1388_));
 OAI21_X1 _5080_ (.A(_1361_),
    .B1(_1388_),
    .B2(_1384_),
    .ZN(_1389_));
 INV_X1 _5081_ (.A(_1389_),
    .ZN(_1390_));
 NOR2_X1 _5082_ (.A1(_1384_),
    .A2(_1388_),
    .ZN(_1391_));
 XNOR2_X1 _5083_ (.A(_1391_),
    .B(_1361_),
    .ZN(_1392_));
 XNOR2_X1 _5084_ (.A(_1379_),
    .B(_1381_),
    .ZN(_1393_));
 XOR2_X1 _5085_ (.A(_1366_),
    .B(_1367_),
    .Z(_1394_));
 XNOR2_X1 _5086_ (.A(_2336_),
    .B(_1394_),
    .ZN(_1395_));
 NAND2_X1 _5087_ (.A1(_1181_),
    .A2(_1182_),
    .ZN(_1397_));
 XNOR2_X1 _5088_ (.A(_1397_),
    .B(_1184_),
    .ZN(_1398_));
 NAND2_X1 _5089_ (.A1(\iir1.y[0] ),
    .A2(_1398_),
    .ZN(_1399_));
 XNOR2_X1 _5090_ (.A(\iir1.y[1] ),
    .B(_1365_),
    .ZN(_1400_));
 XOR2_X1 _5091_ (.A(_1399_),
    .B(_1400_),
    .Z(_1401_));
 AND2_X1 _5092_ (.A1(\iir1.y[3] ),
    .A2(_1401_),
    .ZN(_1402_));
 NOR2_X1 _5093_ (.A1(_1399_),
    .A2(_1400_),
    .ZN(_1403_));
 OAI21_X1 _5094_ (.A(_1395_),
    .B1(_1402_),
    .B2(_1403_),
    .ZN(_1404_));
 OR3_X1 _5095_ (.A1(_1403_),
    .A2(_1402_),
    .A3(_1395_),
    .ZN(_1405_));
 AND2_X1 _5096_ (.A1(_1404_),
    .A2(_1405_),
    .ZN(_1406_));
 NAND2_X1 _5097_ (.A1(\iir1.y[7] ),
    .A2(_1406_),
    .ZN(_1408_));
 NAND2_X1 _5098_ (.A1(_1404_),
    .A2(_1408_),
    .ZN(_1409_));
 XOR2_X1 _5099_ (.A(_1370_),
    .B(_1372_),
    .Z(_1410_));
 XNOR2_X1 _5100_ (.A(_1410_),
    .B(_1376_),
    .ZN(_1411_));
 XOR2_X1 _5101_ (.A(_1409_),
    .B(_1411_),
    .Z(_1412_));
 NAND2_X1 _5102_ (.A1(\iir1.y[8] ),
    .A2(_1412_),
    .ZN(_1413_));
 NAND2_X1 _5103_ (.A1(_1409_),
    .A2(_1411_),
    .ZN(_1414_));
 AOI21_X1 _5104_ (.A(_1393_),
    .B1(_1413_),
    .B2(_1414_),
    .ZN(_1415_));
 XOR2_X1 _5105_ (.A(_1362_),
    .B(_1387_),
    .Z(_1416_));
 AND2_X1 _5106_ (.A1(_1415_),
    .A2(_1416_),
    .ZN(_1417_));
 XOR2_X1 _5107_ (.A(_1415_),
    .B(_1416_),
    .Z(_1419_));
 XNOR2_X1 _5108_ (.A(\iir1.y[7] ),
    .B(_1406_),
    .ZN(_1420_));
 XOR2_X1 _5109_ (.A(_1181_),
    .B(_1182_),
    .Z(_1421_));
 NAND2_X1 _5110_ (.A1(\iir1.y[1] ),
    .A2(_1421_),
    .ZN(_1422_));
 XNOR2_X1 _5111_ (.A(\iir1.y[0] ),
    .B(_1398_),
    .ZN(_1423_));
 NOR2_X1 _5112_ (.A1(_1422_),
    .A2(_1423_),
    .ZN(_1424_));
 XOR2_X1 _5113_ (.A(_1422_),
    .B(_1423_),
    .Z(_1425_));
 AOI21_X1 _5114_ (.A(_1424_),
    .B1(_1425_),
    .B2(\iir1.y[2] ),
    .ZN(_1426_));
 XNOR2_X1 _5115_ (.A(\iir1.y[3] ),
    .B(_1401_),
    .ZN(_1427_));
 XOR2_X1 _5116_ (.A(_1426_),
    .B(_1427_),
    .Z(_1428_));
 NAND2_X1 _5117_ (.A1(\iir1.y[6] ),
    .A2(_1428_),
    .ZN(_1430_));
 OR2_X1 _5118_ (.A1(_1426_),
    .A2(_1427_),
    .ZN(_1431_));
 AOI21_X1 _5119_ (.A(_1420_),
    .B1(_1430_),
    .B2(_1431_),
    .ZN(_1432_));
 XOR2_X1 _5120_ (.A(\iir1.y[8] ),
    .B(_1412_),
    .Z(_1433_));
 AND3_X1 _5121_ (.A1(_1414_),
    .A2(_1413_),
    .A3(_1393_),
    .ZN(_1434_));
 NOR2_X1 _5122_ (.A1(_1415_),
    .A2(_1434_),
    .ZN(_1435_));
 NAND3_X1 _5123_ (.A1(_1432_),
    .A2(_1433_),
    .A3(_1435_),
    .ZN(_1436_));
 NAND2_X1 _5124_ (.A1(_1432_),
    .A2(_1433_),
    .ZN(_1437_));
 XNOR2_X1 _5125_ (.A(_1437_),
    .B(_1435_),
    .ZN(_1438_));
 INV_X1 _5126_ (.A(_1438_),
    .ZN(_1439_));
 XNOR2_X1 _5127_ (.A(\iir1.y[6] ),
    .B(_1428_),
    .ZN(_1441_));
 XOR2_X1 _5128_ (.A(_1179_),
    .B(_1180_),
    .Z(_1442_));
 XNOR2_X1 _5129_ (.A(\iir1.x2[0] ),
    .B(_1442_),
    .ZN(_1443_));
 XNOR2_X1 _5130_ (.A(\iir1.y[1] ),
    .B(_1421_),
    .ZN(_1444_));
 NOR3_X1 _5131_ (.A1(_0737_),
    .A2(_1443_),
    .A3(_1444_),
    .ZN(_1445_));
 NOR2_X1 _5132_ (.A1(_0737_),
    .A2(_1443_),
    .ZN(_1446_));
 XNOR2_X1 _5133_ (.A(_1446_),
    .B(_1444_),
    .ZN(_1447_));
 AOI21_X1 _5134_ (.A(_1445_),
    .B1(_1447_),
    .B2(\iir1.y[4] ),
    .ZN(_1448_));
 XNOR2_X1 _5135_ (.A(\iir1.y[2] ),
    .B(_1425_),
    .ZN(_1449_));
 XOR2_X1 _5136_ (.A(_1448_),
    .B(_1449_),
    .Z(_1450_));
 NAND2_X1 _5137_ (.A1(\iir1.y[5] ),
    .A2(_1450_),
    .ZN(_1452_));
 OR2_X1 _5138_ (.A1(_1448_),
    .A2(_1449_),
    .ZN(_1453_));
 AOI21_X1 _5139_ (.A(_1441_),
    .B1(_1452_),
    .B2(_1453_),
    .ZN(_1454_));
 AND3_X1 _5140_ (.A1(_1431_),
    .A2(_1430_),
    .A3(_1420_),
    .ZN(_1455_));
 NOR2_X1 _5141_ (.A1(_1432_),
    .A2(_1455_),
    .ZN(_1456_));
 NAND2_X1 _5142_ (.A1(_1454_),
    .A2(_1456_),
    .ZN(_1457_));
 XNOR2_X1 _5143_ (.A(_1432_),
    .B(_1433_),
    .ZN(_1458_));
 NOR2_X1 _5144_ (.A1(_1457_),
    .A2(_1458_),
    .ZN(_1459_));
 XNOR2_X1 _5145_ (.A(_0737_),
    .B(_1443_),
    .ZN(_1460_));
 INV_X1 _5146_ (.A(_1460_),
    .ZN(_1461_));
 NAND2_X1 _5147_ (.A1(\iir1.y[3] ),
    .A2(_1461_),
    .ZN(_1463_));
 XNOR2_X1 _5148_ (.A(\iir1.y[4] ),
    .B(_1447_),
    .ZN(_1464_));
 NOR2_X1 _5149_ (.A1(_1463_),
    .A2(_1464_),
    .ZN(_1465_));
 XNOR2_X1 _5150_ (.A(\iir1.y[5] ),
    .B(_1450_),
    .ZN(_1466_));
 INV_X1 _5151_ (.A(_1466_),
    .ZN(_1467_));
 AND3_X1 _5152_ (.A1(_1453_),
    .A2(_1452_),
    .A3(_1441_),
    .ZN(_1468_));
 NOR2_X1 _5153_ (.A1(_1454_),
    .A2(_1468_),
    .ZN(_1469_));
 NAND3_X1 _5154_ (.A1(_1465_),
    .A2(_1467_),
    .A3(_1469_),
    .ZN(_1470_));
 XNOR2_X1 _5155_ (.A(_1454_),
    .B(_1456_),
    .ZN(_1471_));
 XOR2_X1 _5156_ (.A(_1470_),
    .B(_1471_),
    .Z(_1472_));
 XOR2_X1 _5157_ (.A(\iir1.y[3] ),
    .B(_1460_),
    .Z(_1474_));
 NAND2_X1 _5158_ (.A1(\iir1.y[1] ),
    .A2(\iir1.t1[1] ),
    .ZN(_1475_));
 XNOR2_X1 _5159_ (.A(\iir1.x2[0] ),
    .B(_1178_),
    .ZN(_1476_));
 XOR2_X1 _5160_ (.A(_1475_),
    .B(_1476_),
    .Z(_1477_));
 NAND2_X1 _5161_ (.A1(\iir1.y[2] ),
    .A2(_1477_),
    .ZN(_1478_));
 OR2_X1 _5162_ (.A1(_1475_),
    .A2(_1476_),
    .ZN(_1479_));
 AOI21_X1 _5163_ (.A(_1474_),
    .B1(_1478_),
    .B2(_1479_),
    .ZN(_1480_));
 XOR2_X1 _5164_ (.A(_1463_),
    .B(_1464_),
    .Z(_1481_));
 AND3_X1 _5165_ (.A1(_1467_),
    .A2(_1480_),
    .A3(_1481_),
    .ZN(_1482_));
 NAND2_X1 _5166_ (.A1(_1465_),
    .A2(_1467_),
    .ZN(_1483_));
 XNOR2_X1 _5167_ (.A(_1483_),
    .B(_1469_),
    .ZN(_1485_));
 NAND2_X1 _5168_ (.A1(_1482_),
    .A2(_1485_),
    .ZN(_1486_));
 XOR2_X1 _5169_ (.A(\iir1.y[1] ),
    .B(\iir1.t1[1] ),
    .Z(_1487_));
 NAND3_X1 _5170_ (.A1(\iir1.y[0] ),
    .A2(\iir1.t1[0] ),
    .A3(_1487_),
    .ZN(_1488_));
 XNOR2_X1 _5171_ (.A(\iir1.y[2] ),
    .B(_1477_),
    .ZN(_1489_));
 NOR2_X1 _5172_ (.A1(_1488_),
    .A2(_1489_),
    .ZN(_1490_));
 AND3_X1 _5173_ (.A1(_1479_),
    .A2(_1478_),
    .A3(_1474_),
    .ZN(_1491_));
 NOR2_X1 _5174_ (.A1(_1480_),
    .A2(_1491_),
    .ZN(_1492_));
 NAND2_X1 _5175_ (.A1(_1490_),
    .A2(_1492_),
    .ZN(_1493_));
 XNOR2_X1 _5176_ (.A(_1480_),
    .B(_1481_),
    .ZN(_1494_));
 OR2_X1 _5177_ (.A1(_1493_),
    .A2(_1494_),
    .ZN(_1496_));
 AOI21_X1 _5178_ (.A(_1465_),
    .B1(_1480_),
    .B2(_1481_),
    .ZN(_1497_));
 XNOR2_X1 _5179_ (.A(_1466_),
    .B(_1497_),
    .ZN(_1498_));
 OR2_X1 _5180_ (.A1(_1496_),
    .A2(_1498_),
    .ZN(_1499_));
 XNOR2_X1 _5181_ (.A(_1482_),
    .B(_1485_),
    .ZN(_1500_));
 OAI21_X1 _5182_ (.A(_1486_),
    .B1(_1499_),
    .B2(_1500_),
    .ZN(_1501_));
 NAND2_X1 _5183_ (.A1(_1472_),
    .A2(_1501_),
    .ZN(_1502_));
 OAI21_X1 _5184_ (.A(_1502_),
    .B1(_1471_),
    .B2(_1470_),
    .ZN(_1503_));
 XOR2_X1 _5185_ (.A(_1457_),
    .B(_1458_),
    .Z(_1504_));
 AOI21_X1 _5186_ (.A(_1459_),
    .B1(_1503_),
    .B2(_1504_),
    .ZN(_1505_));
 OAI21_X1 _5187_ (.A(_1436_),
    .B1(_1439_),
    .B2(_1505_),
    .ZN(_1507_));
 AOI21_X1 _5188_ (.A(_1417_),
    .B1(_1419_),
    .B2(_1507_),
    .ZN(_1508_));
 INV_X1 _5189_ (.A(_1508_),
    .ZN(_1509_));
 AOI21_X1 _5190_ (.A(_1390_),
    .B1(_1392_),
    .B2(_1509_),
    .ZN(_1510_));
 OAI21_X1 _5191_ (.A(_1358_),
    .B1(_1359_),
    .B2(_1510_),
    .ZN(_1511_));
 AOI21_X1 _5192_ (.A(_1339_),
    .B1(_1340_),
    .B2(_1511_),
    .ZN(_1512_));
 NOR3_X1 _5193_ (.A1(\iir1.y[9] ),
    .A2(_0005_),
    .A3(_2721_),
    .ZN(_1513_));
 XNOR2_X1 _5194_ (.A(\iir1.y[5] ),
    .B(_1946_),
    .ZN(_1514_));
 NAND2_X1 _5195_ (.A1(_1550_),
    .A2(_1327_),
    .ZN(_1515_));
 OAI21_X1 _5196_ (.A(_1324_),
    .B1(_1326_),
    .B2(_1291_),
    .ZN(_1516_));
 OAI21_X1 _5197_ (.A(_1296_),
    .B1(_1298_),
    .B2(\iir1.x2[9] ),
    .ZN(_1518_));
 AOI22_X1 _5198_ (.A1(_1304_),
    .A2(_1315_),
    .B1(_1316_),
    .B2(_1302_),
    .ZN(_1519_));
 OAI21_X1 _5199_ (.A(\iir1.x2[10] ),
    .B1(\iir1.x2[9] ),
    .B2(\iir1.x[9] ),
    .ZN(_1520_));
 NAND3_X1 _5200_ (.A1(\iir1.x[9] ),
    .A2(\iir1.x2[10] ),
    .A3(\iir1.x2[9] ),
    .ZN(_1521_));
 INV_X1 _5201_ (.A(_1521_),
    .ZN(_1522_));
 NOR2_X1 _5202_ (.A1(_1520_),
    .A2(_1522_),
    .ZN(_1523_));
 AND2_X1 _5203_ (.A1(_1306_),
    .A2(_1313_),
    .ZN(_1524_));
 NOR2_X1 _5204_ (.A1(_1305_),
    .A2(_1314_),
    .ZN(_1525_));
 NOR2_X1 _5205_ (.A1(_1524_),
    .A2(_1525_),
    .ZN(_1526_));
 XNOR2_X1 _5206_ (.A(\iir1.x[10] ),
    .B(\iir1.x2[10] ),
    .ZN(_1527_));
 XNOR2_X1 _5207_ (.A(\iir1.x1[9] ),
    .B(_1307_),
    .ZN(_1529_));
 INV_X1 _5208_ (.A(_1312_),
    .ZN(_1530_));
 AOI21_X1 _5209_ (.A(_1530_),
    .B1(_1307_),
    .B2(\iir1.x1[5] ),
    .ZN(_1531_));
 OR2_X1 _5210_ (.A1(_1309_),
    .A2(_1531_),
    .ZN(_1532_));
 XOR2_X1 _5211_ (.A(_1529_),
    .B(_1532_),
    .Z(_1533_));
 XNOR2_X1 _5212_ (.A(_0010_),
    .B(_1533_),
    .ZN(_1534_));
 XNOR2_X1 _5213_ (.A(_1527_),
    .B(_1534_),
    .ZN(_1535_));
 XNOR2_X1 _5214_ (.A(_1526_),
    .B(_1535_),
    .ZN(_1536_));
 XNOR2_X1 _5215_ (.A(_1523_),
    .B(_1536_),
    .ZN(_1537_));
 XOR2_X1 _5216_ (.A(_1519_),
    .B(_1537_),
    .Z(_1538_));
 XNOR2_X1 _5217_ (.A(_1518_),
    .B(_1538_),
    .ZN(_1540_));
 INV_X1 _5218_ (.A(_1318_),
    .ZN(_1541_));
 NAND2_X1 _5219_ (.A1(_1292_),
    .A2(_1541_),
    .ZN(_1542_));
 OR2_X1 _5220_ (.A1(_1294_),
    .A2(_1317_),
    .ZN(_1543_));
 AOI21_X1 _5221_ (.A(_1540_),
    .B1(_1542_),
    .B2(_1543_),
    .ZN(_1544_));
 AND3_X1 _5222_ (.A1(_1543_),
    .A2(_1542_),
    .A3(_1540_),
    .ZN(_1545_));
 NOR2_X1 _5223_ (.A1(_1544_),
    .A2(_1545_),
    .ZN(_1546_));
 XOR2_X1 _5224_ (.A(_1516_),
    .B(_1546_),
    .Z(_1547_));
 XNOR2_X1 _5225_ (.A(\iir1.y[4] ),
    .B(_1547_),
    .ZN(_1548_));
 XNOR2_X1 _5226_ (.A(_1515_),
    .B(_1548_),
    .ZN(_1549_));
 XNOR2_X1 _5227_ (.A(_1514_),
    .B(_1549_),
    .ZN(_1551_));
 OR2_X1 _5228_ (.A1(_1572_),
    .A2(_1329_),
    .ZN(_1552_));
 NAND2_X1 _5229_ (.A1(_1289_),
    .A2(_1328_),
    .ZN(_1553_));
 AOI21_X1 _5230_ (.A(_1551_),
    .B1(_1552_),
    .B2(_1553_),
    .ZN(_1554_));
 AND3_X1 _5231_ (.A1(_1553_),
    .A2(_1552_),
    .A3(_1551_),
    .ZN(_1555_));
 OR2_X1 _5232_ (.A1(_1554_),
    .A2(_1555_),
    .ZN(_1556_));
 OR2_X1 _5233_ (.A1(_0005_),
    .A2(_2720_),
    .ZN(_1557_));
 AOI21_X1 _5234_ (.A(_1556_),
    .B1(_1557_),
    .B2(_2572_),
    .ZN(_1558_));
 AND3_X1 _5235_ (.A1(_2572_),
    .A2(_1557_),
    .A3(_1556_),
    .ZN(_1559_));
 OR2_X1 _5236_ (.A1(_1558_),
    .A2(_1559_),
    .ZN(_1560_));
 OR2_X1 _5237_ (.A1(_1332_),
    .A2(_1333_),
    .ZN(_1562_));
 NAND2_X1 _5238_ (.A1(_1287_),
    .A2(_1331_),
    .ZN(_1563_));
 AOI21_X1 _5239_ (.A(_1560_),
    .B1(_1562_),
    .B2(_1563_),
    .ZN(_1564_));
 AND3_X1 _5240_ (.A1(_1563_),
    .A2(_1562_),
    .A3(_1560_),
    .ZN(_1565_));
 OR2_X1 _5241_ (.A1(_1564_),
    .A2(_1565_),
    .ZN(_1566_));
 XNOR2_X1 _5242_ (.A(_1513_),
    .B(_1566_),
    .ZN(_1567_));
 XNOR2_X1 _5243_ (.A(_1336_),
    .B(_1567_),
    .ZN(_1568_));
 XOR2_X1 _5244_ (.A(_1512_),
    .B(_1568_),
    .Z(_1569_));
 XNOR2_X1 _5245_ (.A(_0004_),
    .B(_1569_),
    .ZN(_1570_));
 NAND2_X1 _5246_ (.A1(_0914_),
    .A2(_1570_),
    .ZN(_1571_));
 INV_X1 _5247_ (.A(_1569_),
    .ZN(_1573_));
 OAI21_X1 _5248_ (.A(_1571_),
    .B1(_1573_),
    .B2(_0004_),
    .ZN(_1574_));
 NAND2_X1 _5249_ (.A1(_1336_),
    .A2(_1567_),
    .ZN(_1575_));
 OAI21_X1 _5250_ (.A(_1575_),
    .B1(_1568_),
    .B2(_1512_),
    .ZN(_1576_));
 NOR4_X1 _5251_ (.A1(\iir1.y[9] ),
    .A2(_0005_),
    .A3(_2721_),
    .A4(_1566_),
    .ZN(_1577_));
 OR2_X1 _5252_ (.A1(_1564_),
    .A2(_1577_),
    .ZN(_1578_));
 NAND2_X1 _5253_ (.A1(\iir1.y[5] ),
    .A2(_1946_),
    .ZN(_1579_));
 XNOR2_X1 _5254_ (.A(_2720_),
    .B(_1579_),
    .ZN(_1580_));
 AND2_X1 _5255_ (.A1(\iir1.y[4] ),
    .A2(_1547_),
    .ZN(_1581_));
 OAI21_X1 _5256_ (.A(_1535_),
    .B1(_1525_),
    .B2(_1524_),
    .ZN(_1582_));
 NAND2_X1 _5257_ (.A1(_1523_),
    .A2(_1536_),
    .ZN(_1584_));
 NAND2_X1 _5258_ (.A1(_1582_),
    .A2(_1584_),
    .ZN(_1585_));
 NOR2_X1 _5259_ (.A1(\iir1.x[10] ),
    .A2(_1295_),
    .ZN(_1586_));
 INV_X1 _5260_ (.A(_0010_),
    .ZN(_1587_));
 NAND2_X1 _5261_ (.A1(_1587_),
    .A2(_1533_),
    .ZN(_1588_));
 INV_X1 _5262_ (.A(_1534_),
    .ZN(_1589_));
 OAI21_X1 _5263_ (.A(_1588_),
    .B1(_1589_),
    .B2(_1527_),
    .ZN(_1590_));
 NOR2_X1 _5264_ (.A1(_1529_),
    .A2(_1532_),
    .ZN(_1591_));
 INV_X1 _5265_ (.A(net51),
    .ZN(_1592_));
 NOR3_X1 _5266_ (.A1(\iir1.x1[9] ),
    .A2(\iir1.x1[8] ),
    .A3(\iir1.x1[7] ),
    .ZN(_1593_));
 AOI21_X1 _5267_ (.A(_1592_),
    .B1(_1593_),
    .B2(_1233_),
    .ZN(_1595_));
 NOR2_X1 _5268_ (.A1(_1591_),
    .A2(_1595_),
    .ZN(_1596_));
 XNOR2_X1 _5269_ (.A(_0010_),
    .B(_1596_),
    .ZN(_1597_));
 XOR2_X1 _5270_ (.A(_1527_),
    .B(_1597_),
    .Z(_1598_));
 XNOR2_X1 _5271_ (.A(_1590_),
    .B(_1598_),
    .ZN(_1599_));
 XNOR2_X1 _5272_ (.A(_1586_),
    .B(_1599_),
    .ZN(_1600_));
 XNOR2_X1 _5273_ (.A(_1585_),
    .B(_1600_),
    .ZN(_1601_));
 XNOR2_X1 _5274_ (.A(_1522_),
    .B(_1601_),
    .ZN(_1602_));
 AND2_X1 _5275_ (.A1(_1518_),
    .A2(_1538_),
    .ZN(_1603_));
 NOR2_X1 _5276_ (.A1(_1519_),
    .A2(_1537_),
    .ZN(_1604_));
 OAI21_X1 _5277_ (.A(_1602_),
    .B1(_1603_),
    .B2(_1604_),
    .ZN(_1606_));
 OR3_X1 _5278_ (.A1(_1604_),
    .A2(_1603_),
    .A3(_1602_),
    .ZN(_1607_));
 NAND2_X1 _5279_ (.A1(_1606_),
    .A2(_1607_),
    .ZN(_1608_));
 AOI21_X1 _5280_ (.A(_1544_),
    .B1(_1546_),
    .B2(_1516_),
    .ZN(_1609_));
 XOR2_X1 _5281_ (.A(_1608_),
    .B(_1609_),
    .Z(_1610_));
 XOR2_X1 _5282_ (.A(_1581_),
    .B(_1610_),
    .Z(_1611_));
 XOR2_X1 _5283_ (.A(_2279_),
    .B(_1611_),
    .Z(_1612_));
 NOR2_X1 _5284_ (.A1(_1514_),
    .A2(_1549_),
    .ZN(_1613_));
 NOR2_X1 _5285_ (.A1(_1515_),
    .A2(_1548_),
    .ZN(_1614_));
 OAI21_X1 _5286_ (.A(_1612_),
    .B1(_1613_),
    .B2(_1614_),
    .ZN(_1615_));
 OR3_X1 _5287_ (.A1(_1614_),
    .A2(_1613_),
    .A3(_1612_),
    .ZN(_1617_));
 NAND2_X1 _5288_ (.A1(_1615_),
    .A2(_1617_),
    .ZN(_1618_));
 XOR2_X1 _5289_ (.A(_1580_),
    .B(_1618_),
    .Z(_1619_));
 OAI21_X1 _5290_ (.A(_1619_),
    .B1(_1558_),
    .B2(_1554_),
    .ZN(_1620_));
 OR3_X1 _5291_ (.A1(_1554_),
    .A2(_1558_),
    .A3(_1619_),
    .ZN(_1621_));
 AND2_X1 _5292_ (.A1(_1620_),
    .A2(_1621_),
    .ZN(_1622_));
 XOR2_X1 _5293_ (.A(_1578_),
    .B(_1622_),
    .Z(_1623_));
 XOR2_X1 _5294_ (.A(_1576_),
    .B(_1623_),
    .Z(_1624_));
 XNOR2_X1 _5295_ (.A(\iir1.y2[10] ),
    .B(_1624_),
    .ZN(_1625_));
 XNOR2_X1 _5296_ (.A(_1574_),
    .B(_1625_),
    .ZN(_1626_));
 NAND2_X1 _5297_ (.A1(_0913_),
    .A2(_1626_),
    .ZN(_1628_));
 INV_X1 _5298_ (.A(_1574_),
    .ZN(_1629_));
 OAI21_X1 _5299_ (.A(_1628_),
    .B1(_1625_),
    .B2(_1629_),
    .ZN(_1630_));
 NAND2_X1 _5300_ (.A1(\iir1.y2[9] ),
    .A2(\iir1.y2[7] ),
    .ZN(_1631_));
 XNOR2_X1 _5301_ (.A(_2491_),
    .B(_1631_),
    .ZN(_1632_));
 XOR2_X1 _5302_ (.A(\iir1.y2[10] ),
    .B(_0004_),
    .Z(_1633_));
 XNOR2_X1 _5303_ (.A(_1624_),
    .B(_1633_),
    .ZN(_1634_));
 AND2_X1 _5304_ (.A1(_0138_),
    .A2(_1634_),
    .ZN(_1635_));
 NAND2_X1 _5305_ (.A1(_1578_),
    .A2(_1622_),
    .ZN(_1636_));
 NAND2_X1 _5306_ (.A1(_1576_),
    .A2(_1623_),
    .ZN(_1637_));
 NAND2_X1 _5307_ (.A1(_1636_),
    .A2(_1637_),
    .ZN(_1639_));
 OR2_X1 _5308_ (.A1(_2720_),
    .A2(_1579_),
    .ZN(_1640_));
 OAI21_X1 _5309_ (.A(_1615_),
    .B1(_1618_),
    .B2(_1580_),
    .ZN(_1641_));
 NAND4_X1 _5310_ (.A1(_1516_),
    .A2(_1546_),
    .A3(_1606_),
    .A4(_1607_),
    .ZN(_1642_));
 INV_X1 _5311_ (.A(_1606_),
    .ZN(_1643_));
 AOI21_X1 _5312_ (.A(_1643_),
    .B1(_1607_),
    .B2(_1544_),
    .ZN(_1644_));
 NAND2_X1 _5313_ (.A1(_1585_),
    .A2(_1600_),
    .ZN(_1645_));
 OAI21_X1 _5314_ (.A(_1645_),
    .B1(_1601_),
    .B2(_1521_),
    .ZN(_1646_));
 NAND2_X1 _5315_ (.A1(\iir1.x[10] ),
    .A2(\iir1.x2[10] ),
    .ZN(_1647_));
 NAND2_X1 _5316_ (.A1(_1590_),
    .A2(_1598_),
    .ZN(_1648_));
 INV_X1 _5317_ (.A(_1586_),
    .ZN(_1650_));
 OAI21_X1 _5318_ (.A(_1648_),
    .B1(_1599_),
    .B2(_1650_),
    .ZN(_1651_));
 XNOR2_X1 _5319_ (.A(\iir1.x1[10] ),
    .B(_0010_),
    .ZN(_1652_));
 XNOR2_X1 _5320_ (.A(_1527_),
    .B(_1652_),
    .ZN(_1653_));
 NOR2_X1 _5321_ (.A1(_1527_),
    .A2(_1597_),
    .ZN(_1654_));
 NOR2_X1 _5322_ (.A1(_0010_),
    .A2(_1596_),
    .ZN(_1655_));
 OAI21_X1 _5323_ (.A(_1653_),
    .B1(_1654_),
    .B2(_1655_),
    .ZN(_1656_));
 OR3_X1 _5324_ (.A1(_1655_),
    .A2(_1654_),
    .A3(_1653_),
    .ZN(_1657_));
 AND2_X1 _5325_ (.A1(_1656_),
    .A2(_1657_),
    .ZN(_1658_));
 XNOR2_X1 _5326_ (.A(_1650_),
    .B(_1658_),
    .ZN(_1659_));
 XNOR2_X1 _5327_ (.A(_1651_),
    .B(_1659_),
    .ZN(_1661_));
 XOR2_X1 _5328_ (.A(_1647_),
    .B(_1661_),
    .Z(_1662_));
 XNOR2_X1 _5329_ (.A(_1646_),
    .B(_1662_),
    .ZN(_1663_));
 AND3_X1 _5330_ (.A1(_1642_),
    .A2(_1644_),
    .A3(_1663_),
    .ZN(_1664_));
 AOI21_X1 _5331_ (.A(_1663_),
    .B1(_1644_),
    .B2(_1642_),
    .ZN(_1665_));
 OR2_X1 _5332_ (.A1(_1664_),
    .A2(_1665_),
    .ZN(_1666_));
 NAND2_X1 _5333_ (.A1(\iir1.y[6] ),
    .A2(\iir1.y[5] ),
    .ZN(_1667_));
 XNOR2_X1 _5334_ (.A(_1667_),
    .B(_2333_),
    .ZN(_1668_));
 XOR2_X1 _5335_ (.A(_1666_),
    .B(_1668_),
    .Z(_1669_));
 NAND2_X1 _5336_ (.A1(_2279_),
    .A2(_1611_),
    .ZN(_1670_));
 NAND2_X1 _5337_ (.A1(_1581_),
    .A2(_1610_),
    .ZN(_1672_));
 AOI21_X1 _5338_ (.A(_1669_),
    .B1(_1670_),
    .B2(_1672_),
    .ZN(_1673_));
 AND3_X1 _5339_ (.A1(_1672_),
    .A2(_1670_),
    .A3(_1669_),
    .ZN(_1674_));
 OR2_X1 _5340_ (.A1(_1673_),
    .A2(_1674_),
    .ZN(_1675_));
 XOR2_X1 _5341_ (.A(\iir1.y[10] ),
    .B(_1675_),
    .Z(_1676_));
 XOR2_X1 _5342_ (.A(_1641_),
    .B(_1676_),
    .Z(_1677_));
 XNOR2_X1 _5343_ (.A(_1640_),
    .B(_1677_),
    .ZN(_1678_));
 XOR2_X1 _5344_ (.A(_1620_),
    .B(_1678_),
    .Z(_1679_));
 XNOR2_X1 _5345_ (.A(_1639_),
    .B(_1679_),
    .ZN(_1680_));
 XNOR2_X1 _5346_ (.A(\iir1.y2[10] ),
    .B(_1680_),
    .ZN(_1681_));
 XNOR2_X1 _5347_ (.A(_1635_),
    .B(_1681_),
    .ZN(_1683_));
 XNOR2_X1 _5348_ (.A(_1632_),
    .B(_1683_),
    .ZN(_1684_));
 INV_X1 _5349_ (.A(_1684_),
    .ZN(_1685_));
 NAND2_X1 _5350_ (.A1(_1630_),
    .A2(_1685_),
    .ZN(_1686_));
 XNOR2_X1 _5351_ (.A(_0003_),
    .B(_0911_),
    .ZN(_1687_));
 XOR2_X1 _5352_ (.A(_1630_),
    .B(_1684_),
    .Z(_1688_));
 OAI21_X1 _5353_ (.A(_1686_),
    .B1(_1687_),
    .B2(_1688_),
    .ZN(_1689_));
 MUX2_X1 _5354_ (.A(_0004_),
    .B(_1631_),
    .S(\iir1.y2[8] ),
    .Z(_1690_));
 XNOR2_X1 _5355_ (.A(_0001_),
    .B(_1690_),
    .ZN(_1691_));
 INV_X1 _5356_ (.A(_1691_),
    .ZN(_1692_));
 NAND2_X1 _5357_ (.A1(_1635_),
    .A2(_1681_),
    .ZN(_1694_));
 OAI21_X1 _5358_ (.A(_1694_),
    .B1(_1683_),
    .B2(_1632_),
    .ZN(_1695_));
 INV_X1 _5359_ (.A(_1695_),
    .ZN(_1696_));
 NAND2_X1 _5360_ (.A1(\iir1.y2[8] ),
    .A2(\iir1.y2[10] ),
    .ZN(_1697_));
 XNOR2_X1 _5361_ (.A(_2561_),
    .B(_1697_),
    .ZN(_1698_));
 XNOR2_X1 _5362_ (.A(_1633_),
    .B(_1680_),
    .ZN(_1699_));
 NOR2_X1 _5363_ (.A1(_0004_),
    .A2(_1699_),
    .ZN(_1700_));
 NOR2_X1 _5364_ (.A1(_1620_),
    .A2(_1678_),
    .ZN(_1701_));
 AOI21_X1 _5365_ (.A(_1701_),
    .B1(_1679_),
    .B2(_1639_),
    .ZN(_1702_));
 INV_X1 _5366_ (.A(_1676_),
    .ZN(_1703_));
 NAND2_X1 _5367_ (.A1(_1641_),
    .A2(_1703_),
    .ZN(_1705_));
 OAI21_X1 _5368_ (.A(_1705_),
    .B1(_1677_),
    .B2(_1640_),
    .ZN(_1706_));
 INV_X1 _5369_ (.A(_1675_),
    .ZN(_1707_));
 AOI21_X1 _5370_ (.A(_1673_),
    .B1(_1707_),
    .B2(\iir1.y[10] ),
    .ZN(_1708_));
 NOR2_X1 _5371_ (.A1(\iir1.y[7] ),
    .A2(_1667_),
    .ZN(_1709_));
 XOR2_X1 _5372_ (.A(_1272_),
    .B(_1709_),
    .Z(_1710_));
 INV_X1 _5373_ (.A(_1666_),
    .ZN(_1711_));
 NAND2_X1 _5374_ (.A1(_1711_),
    .A2(_1668_),
    .ZN(_1712_));
 NOR2_X1 _5375_ (.A1(_1286_),
    .A2(\iir1.y[6] ),
    .ZN(_1713_));
 AOI21_X1 _5376_ (.A(_1665_),
    .B1(_1662_),
    .B2(_1646_),
    .ZN(_1714_));
 NAND2_X1 _5377_ (.A1(_1586_),
    .A2(_1658_),
    .ZN(_1716_));
 NAND2_X1 _5378_ (.A1(_1656_),
    .A2(_1716_),
    .ZN(_1717_));
 AOI21_X1 _5379_ (.A(_1650_),
    .B1(_1587_),
    .B2(\iir1.x1[10] ),
    .ZN(_1718_));
 NAND2_X1 _5380_ (.A1(\iir1.x[10] ),
    .A2(_1295_),
    .ZN(_1719_));
 NOR3_X1 _5381_ (.A1(_1592_),
    .A2(_0010_),
    .A3(_1719_),
    .ZN(_1720_));
 NOR2_X1 _5382_ (.A1(\iir1.x1[10] ),
    .A2(_1587_),
    .ZN(_1721_));
 AOI211_X1 _5383_ (.A(_1718_),
    .B(_1720_),
    .C1(_1527_),
    .C2(_1721_),
    .ZN(_1722_));
 XNOR2_X1 _5384_ (.A(_1717_),
    .B(_1722_),
    .ZN(_1723_));
 XOR2_X1 _5385_ (.A(_1647_),
    .B(_1723_),
    .Z(_1724_));
 NOR2_X1 _5386_ (.A1(_1647_),
    .A2(_1661_),
    .ZN(_1725_));
 AND2_X1 _5387_ (.A1(_1651_),
    .A2(_1659_),
    .ZN(_1727_));
 OAI21_X1 _5388_ (.A(_1724_),
    .B1(_1725_),
    .B2(_1727_),
    .ZN(_1728_));
 OR3_X1 _5389_ (.A1(_1727_),
    .A2(_1725_),
    .A3(_1724_),
    .ZN(_1729_));
 AND3_X1 _5390_ (.A1(_1714_),
    .A2(_1728_),
    .A3(_1729_),
    .ZN(_1730_));
 XNOR2_X1 _5391_ (.A(_1713_),
    .B(_1730_),
    .ZN(_1731_));
 XOR2_X1 _5392_ (.A(_1712_),
    .B(_1731_),
    .Z(_1732_));
 XNOR2_X1 _5393_ (.A(_1710_),
    .B(_1732_),
    .ZN(_1733_));
 XOR2_X1 _5394_ (.A(_1708_),
    .B(_1733_),
    .Z(_1734_));
 XNOR2_X1 _5395_ (.A(_1706_),
    .B(_1734_),
    .ZN(_1735_));
 XOR2_X1 _5396_ (.A(_1702_),
    .B(_1735_),
    .Z(_1736_));
 XNOR2_X1 _5397_ (.A(\iir1.y2[10] ),
    .B(_1736_),
    .ZN(_1738_));
 XOR2_X1 _5398_ (.A(_1700_),
    .B(_1738_),
    .Z(_1739_));
 XNOR2_X1 _5399_ (.A(_1698_),
    .B(_1739_),
    .ZN(_1740_));
 XNOR2_X1 _5400_ (.A(_1696_),
    .B(_1740_),
    .ZN(_1741_));
 XNOR2_X1 _5401_ (.A(_1692_),
    .B(_1741_),
    .ZN(_1742_));
 XNOR2_X1 _5402_ (.A(_1689_),
    .B(_1742_),
    .ZN(_1743_));
 NAND3_X1 _5403_ (.A1(_0003_),
    .A2(_0911_),
    .A3(_1743_),
    .ZN(_1744_));
 INV_X1 _5404_ (.A(_1689_),
    .ZN(_1745_));
 OAI21_X1 _5405_ (.A(_1744_),
    .B1(_1742_),
    .B2(_1745_),
    .ZN(_1746_));
 INV_X1 _5406_ (.A(_0001_),
    .ZN(_1747_));
 NOR2_X1 _5407_ (.A1(_1747_),
    .A2(_1690_),
    .ZN(_1749_));
 OAI22_X1 _5408_ (.A1(_1696_),
    .A2(_1740_),
    .B1(_1741_),
    .B2(_1692_),
    .ZN(_1750_));
 MUX2_X1 _5409_ (.A(_0004_),
    .B(_1697_),
    .S(\iir1.y2[9] ),
    .Z(_1751_));
 XOR2_X1 _5410_ (.A(_0008_),
    .B(_1751_),
    .Z(_1752_));
 NOR2_X1 _5411_ (.A1(_1698_),
    .A2(_1739_),
    .ZN(_1753_));
 INV_X1 _5412_ (.A(_1738_),
    .ZN(_1754_));
 AOI21_X1 _5413_ (.A(_1753_),
    .B1(_1754_),
    .B2(_1700_),
    .ZN(_1755_));
 NOR2_X1 _5414_ (.A1(\iir1.y2[9] ),
    .A2(_2704_),
    .ZN(_1756_));
 XNOR2_X1 _5415_ (.A(_1633_),
    .B(_1736_),
    .ZN(_1757_));
 NOR2_X1 _5416_ (.A1(_0004_),
    .A2(_1757_),
    .ZN(_1758_));
 AND2_X1 _5417_ (.A1(_1706_),
    .A2(_1734_),
    .ZN(_1760_));
 NOR2_X1 _5418_ (.A1(_1702_),
    .A2(_1735_),
    .ZN(_1761_));
 NOR2_X1 _5419_ (.A1(_1708_),
    .A2(_1733_),
    .ZN(_1762_));
 AND2_X1 _5420_ (.A1(_1272_),
    .A2(_1709_),
    .ZN(_1763_));
 NOR2_X1 _5421_ (.A1(_1712_),
    .A2(_1731_),
    .ZN(_1764_));
 AOI21_X1 _5422_ (.A(_1764_),
    .B1(_1732_),
    .B2(_1710_),
    .ZN(_1765_));
 INV_X1 _5423_ (.A(_2572_),
    .ZN(_1766_));
 NOR2_X1 _5424_ (.A1(\iir1.y[8] ),
    .A2(_1766_),
    .ZN(_1767_));
 NOR2_X1 _5425_ (.A1(_2574_),
    .A2(_1767_),
    .ZN(_1768_));
 XNOR2_X1 _5426_ (.A(_2442_),
    .B(_1768_),
    .ZN(_1769_));
 INV_X1 _5427_ (.A(_1769_),
    .ZN(_1771_));
 AND2_X1 _5428_ (.A1(_1713_),
    .A2(_1730_),
    .ZN(_1772_));
 NAND2_X1 _5429_ (.A1(_1714_),
    .A2(_1728_),
    .ZN(_1773_));
 NAND2_X1 _5430_ (.A1(_1717_),
    .A2(_1722_),
    .ZN(_1774_));
 OAI21_X1 _5431_ (.A(_1774_),
    .B1(_1723_),
    .B2(_1647_),
    .ZN(_1775_));
 OAI211_X1 _5432_ (.A(\iir1.x1[10] ),
    .B(_1719_),
    .C1(_1586_),
    .C2(_0010_),
    .ZN(_1776_));
 NAND2_X1 _5433_ (.A1(_0010_),
    .A2(_1586_),
    .ZN(_1777_));
 OAI211_X1 _5434_ (.A(_1776_),
    .B(_1777_),
    .C1(_0010_),
    .C2(_1719_),
    .ZN(_1778_));
 XNOR2_X1 _5435_ (.A(_1775_),
    .B(_1778_),
    .ZN(_1779_));
 XNOR2_X1 _5436_ (.A(_1773_),
    .B(_1779_),
    .ZN(_1780_));
 XNOR2_X1 _5437_ (.A(_1772_),
    .B(_1780_),
    .ZN(_1782_));
 XNOR2_X1 _5438_ (.A(_1771_),
    .B(_1782_),
    .ZN(_1783_));
 XOR2_X1 _5439_ (.A(_1765_),
    .B(_1783_),
    .Z(_1784_));
 XOR2_X1 _5440_ (.A(_1763_),
    .B(_1784_),
    .Z(_1785_));
 XOR2_X1 _5441_ (.A(_1762_),
    .B(_1785_),
    .Z(_1786_));
 OR3_X1 _5442_ (.A1(_1760_),
    .A2(_1761_),
    .A3(_1786_),
    .ZN(_1787_));
 OAI21_X1 _5443_ (.A(_1786_),
    .B1(_1761_),
    .B2(_1760_),
    .ZN(_1788_));
 AND2_X1 _5444_ (.A1(_1787_),
    .A2(_1788_),
    .ZN(_1789_));
 XNOR2_X1 _5445_ (.A(_1633_),
    .B(_1789_),
    .ZN(_1790_));
 XNOR2_X1 _5446_ (.A(_1758_),
    .B(_1790_),
    .ZN(_1791_));
 XNOR2_X1 _5447_ (.A(_1756_),
    .B(_1791_),
    .ZN(_1793_));
 XOR2_X1 _5448_ (.A(_1755_),
    .B(_1793_),
    .Z(_1794_));
 XOR2_X1 _5449_ (.A(_1752_),
    .B(_1794_),
    .Z(_1795_));
 XNOR2_X1 _5450_ (.A(_1750_),
    .B(_1795_),
    .ZN(_1796_));
 XNOR2_X1 _5451_ (.A(_1749_),
    .B(_1796_),
    .ZN(_1797_));
 XNOR2_X1 _5452_ (.A(_1746_),
    .B(_1797_),
    .ZN(_1798_));
 XOR2_X1 _5453_ (.A(\iir1.y2[8] ),
    .B(\iir1.y2[6] ),
    .Z(_1799_));
 XNOR2_X1 _5454_ (.A(_1697_),
    .B(_1799_),
    .ZN(_1800_));
 NAND3_X1 _5455_ (.A1(\iir1.y2[7] ),
    .A2(\iir1.y2[5] ),
    .A3(_1800_),
    .ZN(_1801_));
 OAI21_X1 _5456_ (.A(_1801_),
    .B1(_1697_),
    .B2(\iir1.y2[6] ),
    .ZN(_1802_));
 AND2_X1 _5457_ (.A1(_0009_),
    .A2(_1802_),
    .ZN(_1804_));
 XNOR2_X1 _5458_ (.A(_0913_),
    .B(_1626_),
    .ZN(_1805_));
 NAND2_X1 _5459_ (.A1(\iir1.y2[7] ),
    .A2(\iir1.y2[5] ),
    .ZN(_1806_));
 XOR2_X1 _5460_ (.A(_1806_),
    .B(_1800_),
    .Z(_1807_));
 NAND2_X1 _5461_ (.A1(_2491_),
    .A2(_2704_),
    .ZN(_1808_));
 XNOR2_X1 _5462_ (.A(_1340_),
    .B(_1511_),
    .ZN(_1809_));
 XNOR2_X1 _5463_ (.A(_0138_),
    .B(_1809_),
    .ZN(_1810_));
 NAND3_X1 _5464_ (.A1(_1697_),
    .A2(_1808_),
    .A3(_1810_),
    .ZN(_1811_));
 OAI21_X1 _5465_ (.A(_1811_),
    .B1(_1809_),
    .B2(_0004_),
    .ZN(_1812_));
 XOR2_X1 _5466_ (.A(_0914_),
    .B(_1570_),
    .Z(_1813_));
 XNOR2_X1 _5467_ (.A(_1812_),
    .B(_1813_),
    .ZN(_1815_));
 OR2_X1 _5468_ (.A1(_1807_),
    .A2(_1815_),
    .ZN(_1816_));
 NAND2_X1 _5469_ (.A1(_1812_),
    .A2(_1813_),
    .ZN(_1817_));
 AOI21_X1 _5470_ (.A(_1805_),
    .B1(_1816_),
    .B2(_1817_),
    .ZN(_1818_));
 XNOR2_X1 _5471_ (.A(_0009_),
    .B(_1802_),
    .ZN(_1819_));
 AND3_X1 _5472_ (.A1(_1817_),
    .A2(_1816_),
    .A3(_1805_),
    .ZN(_1820_));
 OR2_X1 _5473_ (.A1(_1818_),
    .A2(_1820_),
    .ZN(_1821_));
 NOR2_X1 _5474_ (.A1(_1819_),
    .A2(_1821_),
    .ZN(_1822_));
 NOR2_X1 _5475_ (.A1(_1818_),
    .A2(_1822_),
    .ZN(_1823_));
 XNOR2_X1 _5476_ (.A(_1687_),
    .B(_1688_),
    .ZN(_1824_));
 XOR2_X1 _5477_ (.A(_1823_),
    .B(_1824_),
    .Z(_1826_));
 NAND2_X1 _5478_ (.A1(_1804_),
    .A2(_1826_),
    .ZN(_1827_));
 OAI21_X1 _5479_ (.A(_1827_),
    .B1(_1824_),
    .B2(_1823_),
    .ZN(_1828_));
 NAND2_X1 _5480_ (.A1(_0003_),
    .A2(_0911_),
    .ZN(_1829_));
 XNOR2_X1 _5481_ (.A(_1829_),
    .B(_1743_),
    .ZN(_1830_));
 NAND2_X1 _5482_ (.A1(_1828_),
    .A2(_1830_),
    .ZN(_1831_));
 XOR2_X1 _5483_ (.A(_1828_),
    .B(_1830_),
    .Z(_1832_));
 NAND2_X1 _5484_ (.A1(\iir1.y2[6] ),
    .A2(\iir1.y2[4] ),
    .ZN(_1833_));
 XOR2_X1 _5485_ (.A(\iir1.y2[7] ),
    .B(\iir1.y2[5] ),
    .Z(_1834_));
 XNOR2_X1 _5486_ (.A(_1631_),
    .B(_1834_),
    .ZN(_1835_));
 XOR2_X1 _5487_ (.A(_1833_),
    .B(_1835_),
    .Z(_1837_));
 XNOR2_X1 _5488_ (.A(_1392_),
    .B(_1508_),
    .ZN(_1838_));
 XNOR2_X1 _5489_ (.A(_2704_),
    .B(_1838_),
    .ZN(_1839_));
 AOI22_X1 _5490_ (.A1(_0138_),
    .A2(_1838_),
    .B1(_1839_),
    .B2(\iir1.y2[9] ),
    .ZN(_1840_));
 XOR2_X1 _5491_ (.A(_1510_),
    .B(_1359_),
    .Z(_1841_));
 XNOR2_X1 _5492_ (.A(_1840_),
    .B(_1841_),
    .ZN(_1842_));
 NAND2_X1 _5493_ (.A1(_0908_),
    .A2(_1842_),
    .ZN(_1843_));
 INV_X1 _5494_ (.A(_1841_),
    .ZN(_1844_));
 OAI21_X1 _5495_ (.A(_1843_),
    .B1(_1844_),
    .B2(_1840_),
    .ZN(_1845_));
 NAND2_X1 _5496_ (.A1(_1697_),
    .A2(_1808_),
    .ZN(_1846_));
 XNOR2_X1 _5497_ (.A(_1846_),
    .B(_1810_),
    .ZN(_1848_));
 XNOR2_X1 _5498_ (.A(_1845_),
    .B(_1848_),
    .ZN(_1849_));
 NOR2_X1 _5499_ (.A1(_1837_),
    .A2(_1849_),
    .ZN(_1850_));
 AOI21_X1 _5500_ (.A(_1850_),
    .B1(_1848_),
    .B2(_1845_),
    .ZN(_1851_));
 XNOR2_X1 _5501_ (.A(_1807_),
    .B(_1815_),
    .ZN(_1852_));
 NOR2_X1 _5502_ (.A1(_1851_),
    .A2(_1852_),
    .ZN(_1853_));
 INV_X1 _5503_ (.A(_1835_),
    .ZN(_1854_));
 OAI22_X1 _5504_ (.A1(\iir1.y2[5] ),
    .A2(_1631_),
    .B1(_1833_),
    .B2(_1854_),
    .ZN(_1855_));
 XOR2_X1 _5505_ (.A(_0011_),
    .B(_1855_),
    .Z(_1856_));
 XOR2_X1 _5506_ (.A(_1851_),
    .B(_1852_),
    .Z(_1857_));
 AOI21_X1 _5507_ (.A(_1853_),
    .B1(_1856_),
    .B2(_1857_),
    .ZN(_1859_));
 XNOR2_X1 _5508_ (.A(_1819_),
    .B(_1821_),
    .ZN(_1860_));
 NOR2_X1 _5509_ (.A1(_1859_),
    .A2(_1860_),
    .ZN(_1861_));
 XOR2_X1 _5510_ (.A(_1859_),
    .B(_1860_),
    .Z(_1862_));
 AND2_X1 _5511_ (.A1(_0011_),
    .A2(_1855_),
    .ZN(_1863_));
 AOI21_X1 _5512_ (.A(_1861_),
    .B1(_1862_),
    .B2(_1863_),
    .ZN(_1864_));
 XNOR2_X1 _5513_ (.A(_1804_),
    .B(_1826_),
    .ZN(_1865_));
 XNOR2_X1 _5514_ (.A(_1864_),
    .B(_1865_),
    .ZN(_1866_));
 XOR2_X1 _5515_ (.A(_1863_),
    .B(_1862_),
    .Z(_1867_));
 NAND2_X1 _5516_ (.A1(\iir1.y2[5] ),
    .A2(\iir1.y2[3] ),
    .ZN(_1868_));
 XNOR2_X1 _5517_ (.A(\iir1.y2[6] ),
    .B(\iir1.y2[4] ),
    .ZN(_1870_));
 XOR2_X1 _5518_ (.A(_0912_),
    .B(_1870_),
    .Z(_1871_));
 INV_X1 _5519_ (.A(_1871_),
    .ZN(_1872_));
 OAI22_X1 _5520_ (.A1(\iir1.y2[4] ),
    .A2(_0912_),
    .B1(_1868_),
    .B2(_1872_),
    .ZN(_1873_));
 NAND2_X1 _5521_ (.A1(_0012_),
    .A2(_1873_),
    .ZN(_1874_));
 XOR2_X1 _5522_ (.A(_0908_),
    .B(_1842_),
    .Z(_1875_));
 XNOR2_X1 _5523_ (.A(_1419_),
    .B(_1507_),
    .ZN(_1876_));
 AND2_X1 _5524_ (.A1(_2561_),
    .A2(_1876_),
    .ZN(_1877_));
 XNOR2_X1 _5525_ (.A(\iir1.y2[9] ),
    .B(_1839_),
    .ZN(_1878_));
 XOR2_X1 _5526_ (.A(_1877_),
    .B(_1878_),
    .Z(_1879_));
 AND2_X1 _5527_ (.A1(_1799_),
    .A2(_1879_),
    .ZN(_1881_));
 NOR2_X1 _5528_ (.A1(_1877_),
    .A2(_1878_),
    .ZN(_1882_));
 OAI21_X1 _5529_ (.A(_1875_),
    .B1(_1881_),
    .B2(_1882_),
    .ZN(_1883_));
 XNOR2_X1 _5530_ (.A(_1868_),
    .B(_1871_),
    .ZN(_1884_));
 OR3_X1 _5531_ (.A1(_1882_),
    .A2(_1881_),
    .A3(_1875_),
    .ZN(_1885_));
 AND2_X1 _5532_ (.A1(_1883_),
    .A2(_1885_),
    .ZN(_1886_));
 NAND2_X1 _5533_ (.A1(_1884_),
    .A2(_1886_),
    .ZN(_1887_));
 NAND2_X1 _5534_ (.A1(_1883_),
    .A2(_1887_),
    .ZN(_1888_));
 XNOR2_X1 _5535_ (.A(_1837_),
    .B(_1849_),
    .ZN(_1889_));
 INV_X1 _5536_ (.A(_1889_),
    .ZN(_1890_));
 XOR2_X1 _5537_ (.A(_0012_),
    .B(_1873_),
    .Z(_1892_));
 XNOR2_X1 _5538_ (.A(_1888_),
    .B(_1889_),
    .ZN(_1893_));
 AOI22_X1 _5539_ (.A1(_1888_),
    .A2(_1890_),
    .B1(_1892_),
    .B2(_1893_),
    .ZN(_1894_));
 XNOR2_X1 _5540_ (.A(_1856_),
    .B(_1857_),
    .ZN(_1895_));
 XNOR2_X1 _5541_ (.A(_1894_),
    .B(_1895_),
    .ZN(_1896_));
 NOR2_X1 _5542_ (.A1(_1874_),
    .A2(_1896_),
    .ZN(_1897_));
 NOR2_X1 _5543_ (.A1(_1894_),
    .A2(_1895_),
    .ZN(_1898_));
 OAI21_X1 _5544_ (.A(_1867_),
    .B1(_1897_),
    .B2(_1898_),
    .ZN(_1899_));
 OR3_X1 _5545_ (.A1(_1898_),
    .A2(_1897_),
    .A3(_1867_),
    .ZN(_1900_));
 AND2_X1 _5546_ (.A1(_1899_),
    .A2(_1900_),
    .ZN(_1901_));
 XOR2_X1 _5547_ (.A(_1438_),
    .B(_1505_),
    .Z(_1903_));
 XNOR2_X1 _5548_ (.A(_2491_),
    .B(_1903_),
    .ZN(_1904_));
 OAI22_X1 _5549_ (.A1(_0008_),
    .A2(_1903_),
    .B1(_1904_),
    .B2(_2432_),
    .ZN(_1905_));
 XNOR2_X1 _5550_ (.A(_0030_),
    .B(_1876_),
    .ZN(_1906_));
 NAND2_X1 _5551_ (.A1(_1905_),
    .A2(_1906_),
    .ZN(_1907_));
 XNOR2_X1 _5552_ (.A(\iir1.y2[8] ),
    .B(\iir1.y2[7] ),
    .ZN(_1908_));
 XNOR2_X1 _5553_ (.A(_1905_),
    .B(_1906_),
    .ZN(_1909_));
 OAI21_X1 _5554_ (.A(_1907_),
    .B1(_1908_),
    .B2(_1909_),
    .ZN(_1910_));
 XOR2_X1 _5555_ (.A(_1799_),
    .B(_1879_),
    .Z(_1911_));
 NAND2_X1 _5556_ (.A1(\iir1.y2[5] ),
    .A2(\iir1.y2[4] ),
    .ZN(_1912_));
 NAND2_X1 _5557_ (.A1(\iir1.y2[8] ),
    .A2(\iir1.y2[7] ),
    .ZN(_1914_));
 XOR2_X1 _5558_ (.A(\iir1.y2[5] ),
    .B(\iir1.y2[3] ),
    .Z(_1915_));
 XNOR2_X1 _5559_ (.A(_1914_),
    .B(_1915_),
    .ZN(_1916_));
 XNOR2_X1 _5560_ (.A(_1912_),
    .B(_1916_),
    .ZN(_1917_));
 XOR2_X1 _5561_ (.A(_1910_),
    .B(_1911_),
    .Z(_1918_));
 AOI22_X1 _5562_ (.A1(_1910_),
    .A2(_1911_),
    .B1(_1917_),
    .B2(_1918_),
    .ZN(_1919_));
 XNOR2_X1 _5563_ (.A(_1884_),
    .B(_1886_),
    .ZN(_1920_));
 NOR2_X1 _5564_ (.A1(_1919_),
    .A2(_1920_),
    .ZN(_1921_));
 INV_X1 _5565_ (.A(_0013_),
    .ZN(_1922_));
 NAND3_X1 _5566_ (.A1(\iir1.y2[8] ),
    .A2(\iir1.y2[7] ),
    .A3(_1915_),
    .ZN(_1923_));
 NAND3_X1 _5567_ (.A1(\iir1.y2[5] ),
    .A2(\iir1.y2[4] ),
    .A3(_1916_),
    .ZN(_1925_));
 AND3_X1 _5568_ (.A1(_1922_),
    .A2(_1923_),
    .A3(_1925_),
    .ZN(_1926_));
 AOI21_X1 _5569_ (.A(_1922_),
    .B1(_1923_),
    .B2(_1925_),
    .ZN(_1927_));
 NOR2_X1 _5570_ (.A1(_1926_),
    .A2(_1927_),
    .ZN(_1928_));
 XOR2_X1 _5571_ (.A(_1919_),
    .B(_1920_),
    .Z(_1929_));
 AOI21_X1 _5572_ (.A(_1921_),
    .B1(_1928_),
    .B2(_1929_),
    .ZN(_1930_));
 XNOR2_X1 _5573_ (.A(_1892_),
    .B(_1893_),
    .ZN(_1931_));
 NOR2_X1 _5574_ (.A1(_1930_),
    .A2(_1931_),
    .ZN(_1932_));
 XOR2_X1 _5575_ (.A(_1930_),
    .B(_1931_),
    .Z(_1933_));
 AOI21_X1 _5576_ (.A(_1932_),
    .B1(_1933_),
    .B2(_1927_),
    .ZN(_1934_));
 XNOR2_X1 _5577_ (.A(_1874_),
    .B(_1896_),
    .ZN(_1936_));
 NOR2_X1 _5578_ (.A1(_1934_),
    .A2(_1936_),
    .ZN(_1937_));
 XNOR2_X1 _5579_ (.A(_1934_),
    .B(_1936_),
    .ZN(_1938_));
 XNOR2_X1 _5580_ (.A(_1503_),
    .B(_1504_),
    .ZN(_1939_));
 XNOR2_X1 _5581_ (.A(_2432_),
    .B(_1939_),
    .ZN(_1940_));
 OAI22_X1 _5582_ (.A1(_0001_),
    .A2(_1939_),
    .B1(_1940_),
    .B2(_2430_),
    .ZN(_1941_));
 XNOR2_X1 _5583_ (.A(\iir1.y2[7] ),
    .B(_1904_),
    .ZN(_1942_));
 NAND2_X1 _5584_ (.A1(_1941_),
    .A2(_1942_),
    .ZN(_1943_));
 XNOR2_X1 _5585_ (.A(_1941_),
    .B(_1942_),
    .ZN(_1944_));
 OAI21_X1 _5586_ (.A(_1943_),
    .B1(_1944_),
    .B2(_1870_),
    .ZN(_1945_));
 XOR2_X1 _5587_ (.A(_1908_),
    .B(_1909_),
    .Z(_1947_));
 NAND2_X1 _5588_ (.A1(\iir1.y2[3] ),
    .A2(\iir1.y2[1] ),
    .ZN(_1948_));
 XOR2_X1 _5589_ (.A(\iir1.y2[5] ),
    .B(\iir1.y2[4] ),
    .Z(_1949_));
 XNOR2_X1 _5590_ (.A(_1833_),
    .B(_1949_),
    .ZN(_1950_));
 XNOR2_X1 _5591_ (.A(_1948_),
    .B(_1950_),
    .ZN(_1951_));
 XOR2_X1 _5592_ (.A(_1945_),
    .B(_1947_),
    .Z(_1952_));
 AOI22_X1 _5593_ (.A1(_1945_),
    .A2(_1947_),
    .B1(_1951_),
    .B2(_1952_),
    .ZN(_1953_));
 XNOR2_X1 _5594_ (.A(_1917_),
    .B(_1918_),
    .ZN(_1954_));
 NOR2_X1 _5595_ (.A1(_1953_),
    .A2(_1954_),
    .ZN(_1955_));
 NOR2_X1 _5596_ (.A1(_1506_),
    .A2(\iir1.y2[0] ),
    .ZN(_1956_));
 INV_X1 _5597_ (.A(_0014_),
    .ZN(_1958_));
 NAND3_X1 _5598_ (.A1(\iir1.y2[6] ),
    .A2(_0905_),
    .A3(\iir1.y2[4] ),
    .ZN(_1959_));
 NAND3_X1 _5599_ (.A1(\iir1.y2[3] ),
    .A2(\iir1.y2[1] ),
    .A3(_1950_),
    .ZN(_1960_));
 NAND2_X1 _5600_ (.A1(_1959_),
    .A2(_1960_),
    .ZN(_1961_));
 XNOR2_X1 _5601_ (.A(_1958_),
    .B(_1961_),
    .ZN(_1962_));
 XOR2_X1 _5602_ (.A(_1956_),
    .B(_1962_),
    .Z(_1963_));
 XOR2_X1 _5603_ (.A(_1953_),
    .B(_1954_),
    .Z(_1964_));
 AOI21_X1 _5604_ (.A(_1955_),
    .B1(_1963_),
    .B2(_1964_),
    .ZN(_1965_));
 XNOR2_X1 _5605_ (.A(_1928_),
    .B(_1929_),
    .ZN(_1966_));
 NOR2_X1 _5606_ (.A1(_1965_),
    .A2(_1966_),
    .ZN(_1967_));
 NAND2_X1 _5607_ (.A1(_1956_),
    .A2(_1962_),
    .ZN(_1969_));
 OAI21_X1 _5608_ (.A(_1969_),
    .B1(_1959_),
    .B2(\iir1.y2[1] ),
    .ZN(_1970_));
 XOR2_X1 _5609_ (.A(_1965_),
    .B(_1966_),
    .Z(_1971_));
 AOI21_X1 _5610_ (.A(_1967_),
    .B1(_1970_),
    .B2(_1971_),
    .ZN(_1972_));
 XNOR2_X1 _5611_ (.A(_1927_),
    .B(_1933_),
    .ZN(_1973_));
 OR2_X1 _5612_ (.A1(_1972_),
    .A2(_1973_),
    .ZN(_1974_));
 XOR2_X1 _5613_ (.A(_1972_),
    .B(_1973_),
    .Z(_1975_));
 XOR2_X1 _5614_ (.A(_1963_),
    .B(_1964_),
    .Z(_1976_));
 XNOR2_X1 _5615_ (.A(\iir1.y2[2] ),
    .B(\iir1.y2[0] ),
    .ZN(_1977_));
 XNOR2_X1 _5616_ (.A(\iir1.y2[3] ),
    .B(\iir1.y2[1] ),
    .ZN(_1978_));
 XOR2_X1 _5617_ (.A(_1868_),
    .B(_1978_),
    .Z(_1980_));
 NAND3_X1 _5618_ (.A1(\iir1.y2[2] ),
    .A2(\iir1.y2[0] ),
    .A3(_1980_),
    .ZN(_1981_));
 OAI21_X1 _5619_ (.A(_1981_),
    .B1(_1868_),
    .B2(\iir1.y2[1] ),
    .ZN(_1982_));
 XNOR2_X1 _5620_ (.A(_1977_),
    .B(_1982_),
    .ZN(_1983_));
 XOR2_X1 _5621_ (.A(_1472_),
    .B(_1501_),
    .Z(_1984_));
 INV_X1 _5622_ (.A(_1984_),
    .ZN(_1985_));
 XNOR2_X1 _5623_ (.A(\iir1.y2[6] ),
    .B(_1984_),
    .ZN(_1986_));
 OAI22_X1 _5624_ (.A1(_0003_),
    .A2(_1985_),
    .B1(_1986_),
    .B2(_0905_),
    .ZN(_1987_));
 INV_X1 _5625_ (.A(_1987_),
    .ZN(_1988_));
 XNOR2_X1 _5626_ (.A(_2430_),
    .B(_1940_),
    .ZN(_1989_));
 OR2_X1 _5627_ (.A1(_1988_),
    .A2(_1989_),
    .ZN(_1991_));
 XNOR2_X1 _5628_ (.A(_1988_),
    .B(_1989_),
    .ZN(_1992_));
 INV_X1 _5629_ (.A(_1915_),
    .ZN(_1993_));
 OAI21_X1 _5630_ (.A(_1991_),
    .B1(_1992_),
    .B2(_1993_),
    .ZN(_1994_));
 XOR2_X1 _5631_ (.A(_1870_),
    .B(_1944_),
    .Z(_1995_));
 XOR2_X1 _5632_ (.A(_1994_),
    .B(_1995_),
    .Z(_1996_));
 NAND2_X1 _5633_ (.A1(\iir1.y2[2] ),
    .A2(\iir1.y2[0] ),
    .ZN(_1997_));
 XNOR2_X1 _5634_ (.A(_1997_),
    .B(_1980_),
    .ZN(_1998_));
 AOI22_X1 _5635_ (.A1(_1994_),
    .A2(_1995_),
    .B1(_1996_),
    .B2(_1998_),
    .ZN(_1999_));
 XNOR2_X1 _5636_ (.A(_1951_),
    .B(_1952_),
    .ZN(_2000_));
 XOR2_X1 _5637_ (.A(_1999_),
    .B(_2000_),
    .Z(_2002_));
 INV_X1 _5638_ (.A(_2002_),
    .ZN(_2003_));
 NOR2_X1 _5639_ (.A1(_1983_),
    .A2(_2003_),
    .ZN(_2004_));
 NOR2_X1 _5640_ (.A1(_1999_),
    .A2(_2000_),
    .ZN(_2005_));
 OAI21_X1 _5641_ (.A(_1976_),
    .B1(_2004_),
    .B2(_2005_),
    .ZN(_2006_));
 INV_X1 _5642_ (.A(_2006_),
    .ZN(_2007_));
 NOR2_X1 _5643_ (.A1(_2005_),
    .A2(_2004_),
    .ZN(_2008_));
 XNOR2_X1 _5644_ (.A(_2008_),
    .B(_1976_),
    .ZN(_2009_));
 NAND2_X1 _5645_ (.A1(_1977_),
    .A2(_1982_),
    .ZN(_2010_));
 INV_X1 _5646_ (.A(_2010_),
    .ZN(_2011_));
 AOI21_X1 _5647_ (.A(_2007_),
    .B1(_2009_),
    .B2(_2011_),
    .ZN(_2013_));
 XNOR2_X1 _5648_ (.A(_1970_),
    .B(_1971_),
    .ZN(_2014_));
 OR2_X1 _5649_ (.A1(_2013_),
    .A2(_2014_),
    .ZN(_2015_));
 XOR2_X1 _5650_ (.A(_2013_),
    .B(_2014_),
    .Z(_2016_));
 INV_X1 _5651_ (.A(_2016_),
    .ZN(_2017_));
 XNOR2_X1 _5652_ (.A(_1996_),
    .B(_1998_),
    .ZN(_2018_));
 XNOR2_X1 _5653_ (.A(_1915_),
    .B(_1992_),
    .ZN(_2019_));
 XNOR2_X1 _5654_ (.A(_1499_),
    .B(_1500_),
    .ZN(_2020_));
 XNOR2_X1 _5655_ (.A(_0905_),
    .B(_2020_),
    .ZN(_2021_));
 OAI22_X1 _5656_ (.A1(_0009_),
    .A2(_2020_),
    .B1(_2021_),
    .B2(_2429_),
    .ZN(_2022_));
 INV_X1 _5657_ (.A(_2022_),
    .ZN(_2024_));
 XNOR2_X1 _5658_ (.A(_0905_),
    .B(_1986_),
    .ZN(_2025_));
 XNOR2_X1 _5659_ (.A(_2024_),
    .B(_2025_),
    .ZN(_2026_));
 XNOR2_X1 _5660_ (.A(\iir1.y2[4] ),
    .B(\iir1.y2[2] ),
    .ZN(_2027_));
 NOR2_X1 _5661_ (.A1(_2026_),
    .A2(_2027_),
    .ZN(_2028_));
 NOR2_X1 _5662_ (.A1(_2024_),
    .A2(_2025_),
    .ZN(_2029_));
 OAI21_X1 _5663_ (.A(_2019_),
    .B1(_2028_),
    .B2(_2029_),
    .ZN(_2030_));
 OR3_X1 _5664_ (.A1(_2029_),
    .A2(_2028_),
    .A3(_2019_),
    .ZN(_2031_));
 AND2_X1 _5665_ (.A1(_2030_),
    .A2(_2031_),
    .ZN(_2032_));
 NAND2_X1 _5666_ (.A1(\iir1.y2[4] ),
    .A2(\iir1.y2[2] ),
    .ZN(_2033_));
 XOR2_X1 _5667_ (.A(_1977_),
    .B(_2033_),
    .Z(_2035_));
 NAND2_X1 _5668_ (.A1(_2032_),
    .A2(_2035_),
    .ZN(_2036_));
 AOI21_X1 _5669_ (.A(_2018_),
    .B1(_2036_),
    .B2(_2030_),
    .ZN(_2037_));
 AND3_X1 _5670_ (.A1(_2030_),
    .A2(_2036_),
    .A3(_2018_),
    .ZN(_2038_));
 NOR2_X1 _5671_ (.A1(_2037_),
    .A2(_2038_),
    .ZN(_2039_));
 NOR2_X1 _5672_ (.A1(\iir1.y2[0] ),
    .A2(_2033_),
    .ZN(_2040_));
 AOI21_X1 _5673_ (.A(_2037_),
    .B1(_2039_),
    .B2(_2040_),
    .ZN(_2041_));
 XOR2_X1 _5674_ (.A(_1983_),
    .B(_2002_),
    .Z(_2042_));
 NOR2_X1 _5675_ (.A1(_2041_),
    .A2(_2042_),
    .ZN(_2043_));
 XNOR2_X1 _5676_ (.A(_2010_),
    .B(_2009_),
    .ZN(_2044_));
 XNOR2_X1 _5677_ (.A(_2043_),
    .B(_2044_),
    .ZN(_2046_));
 INV_X1 _5678_ (.A(_2046_),
    .ZN(_2047_));
 XNOR2_X1 _5679_ (.A(_2040_),
    .B(_2039_),
    .ZN(_2048_));
 XNOR2_X1 _5680_ (.A(_1496_),
    .B(_1498_),
    .ZN(_2049_));
 XNOR2_X1 _5681_ (.A(_2429_),
    .B(_2049_),
    .ZN(_2050_));
 OAI22_X1 _5682_ (.A1(_0011_),
    .A2(_2049_),
    .B1(_2050_),
    .B2(_0906_),
    .ZN(_2051_));
 XNOR2_X1 _5683_ (.A(\iir1.y2[4] ),
    .B(_2021_),
    .ZN(_2052_));
 NAND2_X1 _5684_ (.A1(_2051_),
    .A2(_2052_),
    .ZN(_2053_));
 XNOR2_X1 _5685_ (.A(_2051_),
    .B(_2052_),
    .ZN(_2054_));
 OAI21_X1 _5686_ (.A(_2053_),
    .B1(_2054_),
    .B2(_1978_),
    .ZN(_2055_));
 XOR2_X1 _5687_ (.A(_2026_),
    .B(_2027_),
    .Z(_2057_));
 NAND2_X1 _5688_ (.A1(_2055_),
    .A2(_2057_),
    .ZN(_2058_));
 XNOR2_X1 _5689_ (.A(_2055_),
    .B(_2057_),
    .ZN(_2059_));
 NAND2_X1 _5690_ (.A1(_0906_),
    .A2(\iir1.y2[1] ),
    .ZN(_2060_));
 OAI21_X1 _5691_ (.A(_2058_),
    .B1(_2059_),
    .B2(_2060_),
    .ZN(_2061_));
 XNOR2_X1 _5692_ (.A(_2032_),
    .B(_2035_),
    .ZN(_2062_));
 XNOR2_X1 _5693_ (.A(_2061_),
    .B(_2062_),
    .ZN(_2063_));
 NAND3_X1 _5694_ (.A1(\iir1.y2[3] ),
    .A2(\iir1.y2[1] ),
    .A3(_2063_),
    .ZN(_2064_));
 INV_X1 _5695_ (.A(_2062_),
    .ZN(_2065_));
 NAND2_X1 _5696_ (.A1(_2061_),
    .A2(_2065_),
    .ZN(_2066_));
 AOI21_X1 _5697_ (.A(_2048_),
    .B1(_2064_),
    .B2(_2066_),
    .ZN(_2068_));
 XOR2_X1 _5698_ (.A(_2041_),
    .B(_2042_),
    .Z(_2069_));
 NAND2_X1 _5699_ (.A1(_2068_),
    .A2(_2069_),
    .ZN(_2070_));
 NAND2_X1 _5700_ (.A1(_1506_),
    .A2(\iir1.y2[0] ),
    .ZN(_2071_));
 XNOR2_X1 _5701_ (.A(_1493_),
    .B(_1494_),
    .ZN(_2072_));
 XNOR2_X1 _5702_ (.A(_0906_),
    .B(_2072_),
    .ZN(_2073_));
 OAI22_X1 _5703_ (.A1(_0012_),
    .A2(_2072_),
    .B1(_2073_),
    .B2(_1506_),
    .ZN(_2074_));
 XNOR2_X1 _5704_ (.A(\iir1.y2[3] ),
    .B(_2050_),
    .ZN(_2075_));
 NAND2_X1 _5705_ (.A1(_2074_),
    .A2(_2075_),
    .ZN(_2076_));
 XNOR2_X1 _5706_ (.A(_2074_),
    .B(_2075_),
    .ZN(_2077_));
 OAI21_X1 _5707_ (.A(_2076_),
    .B1(_2077_),
    .B2(_1977_),
    .ZN(_2079_));
 XOR2_X1 _5708_ (.A(_1978_),
    .B(_2054_),
    .Z(_2080_));
 XNOR2_X1 _5709_ (.A(_2079_),
    .B(_2080_),
    .ZN(_2081_));
 NOR2_X1 _5710_ (.A1(_2071_),
    .A2(_2081_),
    .ZN(_2082_));
 AOI21_X1 _5711_ (.A(_2082_),
    .B1(_2080_),
    .B2(_2079_),
    .ZN(_2083_));
 XNOR2_X1 _5712_ (.A(_2059_),
    .B(_2060_),
    .ZN(_2084_));
 XNOR2_X1 _5713_ (.A(_2083_),
    .B(_2084_),
    .ZN(_2085_));
 OR2_X1 _5714_ (.A1(_1997_),
    .A2(_2085_),
    .ZN(_2086_));
 OAI21_X1 _5715_ (.A(_2086_),
    .B1(_2084_),
    .B2(_2083_),
    .ZN(_2087_));
 XNOR2_X1 _5716_ (.A(_1948_),
    .B(_2063_),
    .ZN(_2088_));
 XNOR2_X1 _5717_ (.A(_2087_),
    .B(_2088_),
    .ZN(_2090_));
 XNOR2_X1 _5718_ (.A(_1490_),
    .B(_1492_),
    .ZN(_2091_));
 XNOR2_X1 _5719_ (.A(_1506_),
    .B(_2091_),
    .ZN(_2092_));
 OAI22_X1 _5720_ (.A1(_0013_),
    .A2(_2091_),
    .B1(_2092_),
    .B2(_1407_),
    .ZN(_2093_));
 XNOR2_X1 _5721_ (.A(\iir1.y2[2] ),
    .B(_2073_),
    .ZN(_2094_));
 XNOR2_X1 _5722_ (.A(_2093_),
    .B(_2094_),
    .ZN(_2095_));
 XNOR2_X1 _5723_ (.A(_1407_),
    .B(_2095_),
    .ZN(_2096_));
 XOR2_X1 _5724_ (.A(_1488_),
    .B(_1489_),
    .Z(_2097_));
 NAND2_X1 _5725_ (.A1(_1958_),
    .A2(_2097_),
    .ZN(_2098_));
 XNOR2_X1 _5726_ (.A(\iir1.y2[1] ),
    .B(_2097_),
    .ZN(_2099_));
 OAI21_X1 _5727_ (.A(_2098_),
    .B1(_2099_),
    .B2(_2385_),
    .ZN(_2101_));
 XNOR2_X1 _5728_ (.A(\iir1.y2[1] ),
    .B(_2092_),
    .ZN(_2102_));
 XOR2_X1 _5729_ (.A(_2101_),
    .B(_2102_),
    .Z(_2103_));
 NAND2_X1 _5730_ (.A1(\iir1.y2[0] ),
    .A2(_2103_),
    .ZN(_2104_));
 NAND2_X1 _5731_ (.A1(_2101_),
    .A2(_2102_),
    .ZN(_2105_));
 AOI21_X1 _5732_ (.A(_2096_),
    .B1(_2104_),
    .B2(_2105_),
    .ZN(_2106_));
 NAND2_X1 _5733_ (.A1(_2093_),
    .A2(_2094_),
    .ZN(_2107_));
 OAI21_X1 _5734_ (.A(_2107_),
    .B1(_2095_),
    .B2(_1407_),
    .ZN(_2108_));
 XOR2_X1 _5735_ (.A(_1977_),
    .B(_2077_),
    .Z(_2109_));
 XOR2_X1 _5736_ (.A(_2108_),
    .B(_2109_),
    .Z(_2110_));
 AND2_X1 _5737_ (.A1(_2106_),
    .A2(_2110_),
    .ZN(_2112_));
 XOR2_X1 _5738_ (.A(_2071_),
    .B(_2081_),
    .Z(_2113_));
 AND2_X1 _5739_ (.A1(_2112_),
    .A2(_2113_),
    .ZN(_2114_));
 XOR2_X1 _5740_ (.A(_1997_),
    .B(_2085_),
    .Z(_2115_));
 NOR2_X1 _5741_ (.A1(_2114_),
    .A2(_2115_),
    .ZN(_2116_));
 NAND2_X1 _5742_ (.A1(_2114_),
    .A2(_2115_),
    .ZN(_2117_));
 AND2_X1 _5743_ (.A1(_2108_),
    .A2(_2109_),
    .ZN(_2118_));
 XNOR2_X1 _5744_ (.A(_2118_),
    .B(_2113_),
    .ZN(_2119_));
 XNOR2_X1 _5745_ (.A(_2112_),
    .B(_2119_),
    .ZN(_2120_));
 INV_X1 _5746_ (.A(_2110_),
    .ZN(_2121_));
 AOI21_X1 _5747_ (.A(_1487_),
    .B1(\iir1.t1[0] ),
    .B2(\iir1.y[0] ),
    .ZN(_2123_));
 INV_X1 _5748_ (.A(_0015_),
    .ZN(_2124_));
 NAND2_X1 _5749_ (.A1(_2124_),
    .A2(_1488_),
    .ZN(_2125_));
 AOI211_X1 _5750_ (.A(_2123_),
    .B(_2125_),
    .C1(_2385_),
    .C2(_2099_),
    .ZN(_2126_));
 OAI211_X1 _5751_ (.A(_2104_),
    .B(_2126_),
    .C1(_2099_),
    .C2(_2103_),
    .ZN(_2127_));
 AND3_X1 _5752_ (.A1(_2105_),
    .A2(_2104_),
    .A3(_2096_),
    .ZN(_2128_));
 NOR4_X1 _5753_ (.A1(_2106_),
    .A2(_2121_),
    .A3(_2127_),
    .A4(_2128_),
    .ZN(_2129_));
 AOI22_X1 _5754_ (.A1(_2118_),
    .A2(_2113_),
    .B1(_2120_),
    .B2(_2129_),
    .ZN(_2130_));
 AOI211_X1 _5755_ (.A(_2090_),
    .B(_2116_),
    .C1(_2117_),
    .C2(_2130_),
    .ZN(_2131_));
 INV_X1 _5756_ (.A(_2131_),
    .ZN(_2132_));
 AND3_X1 _5757_ (.A1(_2066_),
    .A2(_2064_),
    .A3(_2048_),
    .ZN(_2134_));
 NOR2_X1 _5758_ (.A1(_2068_),
    .A2(_2134_),
    .ZN(_2135_));
 AND2_X1 _5759_ (.A1(_2087_),
    .A2(_2088_),
    .ZN(_2136_));
 XNOR2_X1 _5760_ (.A(_2135_),
    .B(_2136_),
    .ZN(_2137_));
 NOR2_X1 _5761_ (.A1(_2132_),
    .A2(_2137_),
    .ZN(_2138_));
 AOI21_X1 _5762_ (.A(_2138_),
    .B1(_2136_),
    .B2(_2135_),
    .ZN(_2139_));
 XOR2_X1 _5763_ (.A(_2068_),
    .B(_2069_),
    .Z(_2140_));
 INV_X1 _5764_ (.A(_2140_),
    .ZN(_2141_));
 OAI21_X1 _5765_ (.A(_2070_),
    .B1(_2139_),
    .B2(_2141_),
    .ZN(_2142_));
 AOI22_X1 _5766_ (.A1(_2043_),
    .A2(_2044_),
    .B1(_2047_),
    .B2(_2142_),
    .ZN(_2143_));
 OAI21_X1 _5767_ (.A(_2015_),
    .B1(_2017_),
    .B2(_2143_),
    .ZN(_2145_));
 NAND2_X1 _5768_ (.A1(_1975_),
    .A2(_2145_),
    .ZN(_2146_));
 AOI21_X1 _5769_ (.A(_1938_),
    .B1(_1974_),
    .B2(_2146_),
    .ZN(_2147_));
 OAI21_X1 _5770_ (.A(_1901_),
    .B1(_1937_),
    .B2(_2147_),
    .ZN(_2148_));
 AOI21_X1 _5771_ (.A(_1866_),
    .B1(_1899_),
    .B2(_2148_),
    .ZN(_2149_));
 NOR2_X1 _5772_ (.A1(_1864_),
    .A2(_1865_),
    .ZN(_2150_));
 OAI21_X1 _5773_ (.A(_1832_),
    .B1(_2149_),
    .B2(_2150_),
    .ZN(_2151_));
 AOI21_X1 _5774_ (.A(_1798_),
    .B1(_1831_),
    .B2(_2151_),
    .ZN(_2152_));
 AOI21_X1 _5775_ (.A(_2152_),
    .B1(_1797_),
    .B2(_1746_),
    .ZN(_2153_));
 INV_X1 _5776_ (.A(_1751_),
    .ZN(_2154_));
 NAND2_X1 _5777_ (.A1(_0008_),
    .A2(_2154_),
    .ZN(_2156_));
 INV_X1 _5778_ (.A(_1793_),
    .ZN(_2157_));
 OAI22_X1 _5779_ (.A1(_1755_),
    .A2(_2157_),
    .B1(_1794_),
    .B2(_1752_),
    .ZN(_2158_));
 NAND2_X1 _5780_ (.A1(_0138_),
    .A2(_1790_),
    .ZN(_2159_));
 NAND2_X1 _5781_ (.A1(_1762_),
    .A2(_1785_),
    .ZN(_2160_));
 NAND2_X1 _5782_ (.A1(_2160_),
    .A2(_1788_),
    .ZN(_2161_));
 NOR2_X1 _5783_ (.A1(_1765_),
    .A2(_1783_),
    .ZN(_2162_));
 AOI21_X1 _5784_ (.A(_2162_),
    .B1(_1784_),
    .B2(_1763_),
    .ZN(_2163_));
 NOR3_X1 _5785_ (.A1(_2442_),
    .A2(_2574_),
    .A3(_1767_),
    .ZN(_2164_));
 NAND2_X1 _5786_ (.A1(_1772_),
    .A2(_1780_),
    .ZN(_2165_));
 OAI21_X1 _5787_ (.A(_2165_),
    .B1(_1782_),
    .B2(_1771_),
    .ZN(_2167_));
 AOI21_X1 _5788_ (.A(_2647_),
    .B1(_1271_),
    .B2(\iir1.y[9] ),
    .ZN(_2168_));
 NAND2_X1 _5789_ (.A1(_1775_),
    .A2(_1778_),
    .ZN(_2169_));
 OAI211_X1 _5790_ (.A(_1295_),
    .B(_0010_),
    .C1(_1592_),
    .C2(\iir1.x[10] ),
    .ZN(_2170_));
 INV_X1 _5791_ (.A(_1773_),
    .ZN(_2171_));
 OAI211_X1 _5792_ (.A(_2169_),
    .B(_2170_),
    .C1(_1779_),
    .C2(_2171_),
    .ZN(_2172_));
 XOR2_X1 _5793_ (.A(_2168_),
    .B(_2172_),
    .Z(_2173_));
 XOR2_X1 _5794_ (.A(_2167_),
    .B(_2173_),
    .Z(_2174_));
 XOR2_X1 _5795_ (.A(_2164_),
    .B(_2174_),
    .Z(_2175_));
 XNOR2_X1 _5796_ (.A(_2163_),
    .B(_2175_),
    .ZN(_2176_));
 XOR2_X1 _5797_ (.A(_2161_),
    .B(_2176_),
    .Z(_2178_));
 XNOR2_X1 _5798_ (.A(\iir1.y2[10] ),
    .B(_2178_),
    .ZN(_2179_));
 XOR2_X1 _5799_ (.A(_2159_),
    .B(_2179_),
    .Z(_2180_));
 NOR3_X1 _5800_ (.A1(\iir1.y2[9] ),
    .A2(_2704_),
    .A3(_1791_),
    .ZN(_2181_));
 INV_X1 _5801_ (.A(_1757_),
    .ZN(_2182_));
 NOR3_X1 _5802_ (.A1(_0004_),
    .A2(_2182_),
    .A3(_1790_),
    .ZN(_2183_));
 OAI21_X1 _5803_ (.A(_2180_),
    .B1(_2181_),
    .B2(_2183_),
    .ZN(_2184_));
 OR3_X1 _5804_ (.A1(_2183_),
    .A2(_2181_),
    .A3(_2180_),
    .ZN(_2185_));
 AND2_X1 _5805_ (.A1(_2184_),
    .A2(_2185_),
    .ZN(_2186_));
 OAI21_X1 _5806_ (.A(_2186_),
    .B1(\iir1.y2[10] ),
    .B2(_2561_),
    .ZN(_2187_));
 OR3_X1 _5807_ (.A1(_2561_),
    .A2(\iir1.y2[10] ),
    .A3(_2186_),
    .ZN(_2189_));
 AND2_X1 _5808_ (.A1(_2187_),
    .A2(_2189_),
    .ZN(_2190_));
 XOR2_X1 _5809_ (.A(_2158_),
    .B(_2190_),
    .Z(_2191_));
 XNOR2_X1 _5810_ (.A(_2156_),
    .B(_2191_),
    .ZN(_2192_));
 NOR3_X1 _5811_ (.A1(_1747_),
    .A2(_1690_),
    .A3(_1796_),
    .ZN(_2193_));
 AND2_X1 _5812_ (.A1(_1750_),
    .A2(_1795_),
    .ZN(_2194_));
 OAI21_X1 _5813_ (.A(_2192_),
    .B1(_2193_),
    .B2(_2194_),
    .ZN(_2195_));
 OR3_X1 _5814_ (.A1(_2194_),
    .A2(_2193_),
    .A3(_2192_),
    .ZN(_2196_));
 NAND2_X1 _5815_ (.A1(_2195_),
    .A2(_2196_),
    .ZN(_2197_));
 XOR2_X1 _5816_ (.A(_2153_),
    .B(_2197_),
    .Z(_2198_));
 AND3_X1 _5817_ (.A1(_1798_),
    .A2(_1831_),
    .A3(_2151_),
    .ZN(_2200_));
 AND3_X1 _5818_ (.A1(_1866_),
    .A2(_1899_),
    .A3(_2148_),
    .ZN(_2201_));
 NOR2_X1 _5819_ (.A1(_2149_),
    .A2(_2201_),
    .ZN(_2202_));
 OR3_X1 _5820_ (.A1(_1901_),
    .A2(_1937_),
    .A3(_2147_),
    .ZN(_2203_));
 AND2_X1 _5821_ (.A1(_2148_),
    .A2(_2203_),
    .ZN(_2204_));
 AND3_X1 _5822_ (.A1(_1938_),
    .A2(_1974_),
    .A3(_2146_),
    .ZN(_2205_));
 NOR2_X1 _5823_ (.A1(_2147_),
    .A2(_2205_),
    .ZN(_2206_));
 XNOR2_X1 _5824_ (.A(_2016_),
    .B(_2143_),
    .ZN(_2207_));
 XNOR2_X1 _5825_ (.A(_2132_),
    .B(_2137_),
    .ZN(_2208_));
 NOR2_X1 _5826_ (.A1(_2141_),
    .A2(_2208_),
    .ZN(_2209_));
 XNOR2_X1 _5827_ (.A(_2046_),
    .B(_2142_),
    .ZN(_2211_));
 AND2_X1 _5828_ (.A1(_2209_),
    .A2(_2211_),
    .ZN(_2212_));
 AND2_X1 _5829_ (.A1(_2207_),
    .A2(_2212_),
    .ZN(_2213_));
 XOR2_X1 _5830_ (.A(_1975_),
    .B(_2145_),
    .Z(_2214_));
 AND2_X1 _5831_ (.A1(_2213_),
    .A2(_2214_),
    .ZN(_2215_));
 AND2_X1 _5832_ (.A1(_2206_),
    .A2(_2215_),
    .ZN(_2216_));
 AND2_X1 _5833_ (.A1(_2204_),
    .A2(_2216_),
    .ZN(_2217_));
 AND2_X1 _5834_ (.A1(_2202_),
    .A2(_2217_),
    .ZN(_2218_));
 OR3_X1 _5835_ (.A1(_2150_),
    .A2(_2149_),
    .A3(_1832_),
    .ZN(_2219_));
 AND2_X1 _5836_ (.A1(_2151_),
    .A2(_2219_),
    .ZN(_2220_));
 NAND2_X1 _5837_ (.A1(_2218_),
    .A2(_2220_),
    .ZN(_2222_));
 NOR3_X1 _5838_ (.A1(_2152_),
    .A2(_2200_),
    .A3(_2222_),
    .ZN(_2223_));
 OAI21_X1 _5839_ (.A(_1297_),
    .B1(_2198_),
    .B2(_2223_),
    .ZN(_2224_));
 AOI21_X1 _5840_ (.A(_2224_),
    .B1(_2223_),
    .B2(_2198_),
    .ZN(_0086_));
 NOR2_X1 _5841_ (.A1(_2152_),
    .A2(_2200_),
    .ZN(_2225_));
 XOR2_X1 _5842_ (.A(_2225_),
    .B(_2222_),
    .Z(_2226_));
 NOR2_X1 _5843_ (.A1(rst),
    .A2(_2226_),
    .ZN(_0085_));
 OAI21_X1 _5844_ (.A(_1297_),
    .B1(_2218_),
    .B2(_2220_),
    .ZN(_2227_));
 AOI21_X1 _5845_ (.A(_2227_),
    .B1(_2220_),
    .B2(_2218_),
    .ZN(_0084_));
 NOR2_X1 _5846_ (.A1(_2202_),
    .A2(_2217_),
    .ZN(_2228_));
 NOR3_X1 _5847_ (.A1(rst),
    .A2(_2218_),
    .A3(_2228_),
    .ZN(_0083_));
 NOR2_X1 _5848_ (.A1(_2204_),
    .A2(_2216_),
    .ZN(_2230_));
 NOR3_X1 _5849_ (.A1(rst),
    .A2(_2217_),
    .A3(_2230_),
    .ZN(_0082_));
 NOR2_X1 _5850_ (.A1(_2206_),
    .A2(_2215_),
    .ZN(_2231_));
 NOR3_X1 _5851_ (.A1(rst),
    .A2(_2216_),
    .A3(_2231_),
    .ZN(_0081_));
 NOR2_X1 _5852_ (.A1(_2213_),
    .A2(_2214_),
    .ZN(_2232_));
 NOR3_X1 _5853_ (.A1(rst),
    .A2(_2215_),
    .A3(_2232_),
    .ZN(_0080_));
 NOR2_X1 _5854_ (.A1(_2207_),
    .A2(_2212_),
    .ZN(_2233_));
 NOR3_X1 _5855_ (.A1(rst),
    .A2(_2213_),
    .A3(_2233_),
    .ZN(_0079_));
 NOR2_X1 _5856_ (.A1(_2209_),
    .A2(_2211_),
    .ZN(_2234_));
 NOR3_X1 _5857_ (.A1(rst),
    .A2(_2212_),
    .A3(_2234_),
    .ZN(_0078_));
 NAND2_X1 _5858_ (.A1(_2198_),
    .A2(_2223_),
    .ZN(_2236_));
 OAI21_X1 _5859_ (.A(_2195_),
    .B1(_2197_),
    .B2(_2153_),
    .ZN(_2237_));
 NAND2_X1 _5860_ (.A1(_2158_),
    .A2(_2190_),
    .ZN(_2238_));
 NOR2_X1 _5861_ (.A1(_2158_),
    .A2(_2190_),
    .ZN(_2239_));
 OAI21_X1 _5862_ (.A(_2238_),
    .B1(_2239_),
    .B2(_2156_),
    .ZN(_2240_));
 NAND2_X1 _5863_ (.A1(_2184_),
    .A2(_2187_),
    .ZN(_2241_));
 NOR3_X1 _5864_ (.A1(_0004_),
    .A2(_1790_),
    .A3(_2179_),
    .ZN(_2242_));
 NAND3_X1 _5865_ (.A1(\iir1.y2[9] ),
    .A2(\iir1.y2[10] ),
    .A3(_0030_),
    .ZN(_2243_));
 INV_X1 _5866_ (.A(_2175_),
    .ZN(_2244_));
 NOR2_X1 _5867_ (.A1(_2163_),
    .A2(_2244_),
    .ZN(_2246_));
 AOI21_X1 _5868_ (.A(_2246_),
    .B1(_2176_),
    .B2(_2161_),
    .ZN(_2247_));
 AOI22_X1 _5869_ (.A1(_2167_),
    .A2(_2173_),
    .B1(_2174_),
    .B2(_2164_),
    .ZN(_2248_));
 AOI211_X1 _5870_ (.A(_2647_),
    .B(_2172_),
    .C1(_1271_),
    .C2(\iir1.y[9] ),
    .ZN(_2249_));
 XNOR2_X1 _5871_ (.A(_2649_),
    .B(_2249_),
    .ZN(_2250_));
 XNOR2_X1 _5872_ (.A(_2248_),
    .B(_2250_),
    .ZN(_2251_));
 XNOR2_X1 _5873_ (.A(_2247_),
    .B(_2251_),
    .ZN(_2252_));
 XNOR2_X1 _5874_ (.A(_2243_),
    .B(_2252_),
    .ZN(_2253_));
 XNOR2_X1 _5875_ (.A(_2242_),
    .B(_2253_),
    .ZN(_2254_));
 XNOR2_X1 _5876_ (.A(_2241_),
    .B(_2254_),
    .ZN(_2255_));
 XNOR2_X1 _5877_ (.A(_2240_),
    .B(_2255_),
    .ZN(_2257_));
 XNOR2_X1 _5878_ (.A(_2237_),
    .B(_2257_),
    .ZN(_2258_));
 OAI21_X1 _5879_ (.A(_1297_),
    .B1(_2236_),
    .B2(_2258_),
    .ZN(_2259_));
 AOI21_X1 _5880_ (.A(_2259_),
    .B1(_2258_),
    .B2(_2236_),
    .ZN(_0077_));
 XNOR2_X1 _5881_ (.A(_2139_),
    .B(_2141_),
    .ZN(_2260_));
 AND2_X1 _5882_ (.A1(_2208_),
    .A2(_2260_),
    .ZN(_2261_));
 NOR3_X1 _5883_ (.A1(rst),
    .A2(_2209_),
    .A3(_2261_),
    .ZN(_0076_));
 AND2_X1 _5884_ (.A1(_1297_),
    .A2(net59),
    .ZN(_0075_));
 AND2_X1 _5885_ (.A1(_1297_),
    .A2(net83),
    .ZN(_0074_));
 NOR2_X1 _5886_ (.A1(rst),
    .A2(_1286_),
    .ZN(_0073_));
 AND2_X1 _5887_ (.A1(_1297_),
    .A2(net92),
    .ZN(_0072_));
 NOR2_X1 _5888_ (.A1(rst),
    .A2(_2277_),
    .ZN(_0071_));
 AND2_X1 _5889_ (.A1(_1297_),
    .A2(net89),
    .ZN(_0070_));
 AND2_X1 _5890_ (.A1(_1297_),
    .A2(net91),
    .ZN(_0069_));
 AND2_X1 _5891_ (.A1(_1297_),
    .A2(net90),
    .ZN(_0068_));
 AND2_X1 _5892_ (.A1(_1297_),
    .A2(net93),
    .ZN(_0067_));
 AND2_X1 _5893_ (.A1(_1297_),
    .A2(net78),
    .ZN(_0066_));
 NOR2_X1 _5894_ (.A1(rst),
    .A2(_0737_),
    .ZN(_0065_));
 AND2_X1 _5895_ (.A1(_1297_),
    .A2(x[9]),
    .ZN(_0064_));
 AND2_X1 _5896_ (.A1(_1297_),
    .A2(x[8]),
    .ZN(_0063_));
 AND2_X1 _5897_ (.A1(_1297_),
    .A2(x[7]),
    .ZN(_0062_));
 AND2_X1 _5898_ (.A1(_1297_),
    .A2(x[6]),
    .ZN(_0061_));
 AND2_X1 _5899_ (.A1(_1297_),
    .A2(x[5]),
    .ZN(_0060_));
 AND2_X1 _5900_ (.A1(_1297_),
    .A2(x[4]),
    .ZN(_0059_));
 AND2_X1 _5901_ (.A1(_1297_),
    .A2(x[3]),
    .ZN(_0058_));
 AND2_X1 _5902_ (.A1(_1297_),
    .A2(x[2]),
    .ZN(_0057_));
 AND2_X1 _5903_ (.A1(_1297_),
    .A2(x[1]),
    .ZN(_0056_));
 AND2_X1 _5904_ (.A1(_1297_),
    .A2(x[10]),
    .ZN(_0055_));
 AND2_X1 _5905_ (.A1(_1297_),
    .A2(x[0]),
    .ZN(_0054_));
 AND2_X1 _5906_ (.A1(_1297_),
    .A2(net11),
    .ZN(_0053_));
 AND2_X1 _5907_ (.A1(_1297_),
    .A2(net9),
    .ZN(_0052_));
 AND2_X1 _5908_ (.A1(_1297_),
    .A2(net17),
    .ZN(_0051_));
 NOR2_X1 _5909_ (.A1(rst),
    .A2(net2),
    .ZN(_0050_));
 AND2_X1 _5910_ (.A1(_1297_),
    .A2(net37),
    .ZN(_0049_));
 AND2_X1 _5911_ (.A1(_1297_),
    .A2(net4),
    .ZN(_0048_));
 AND2_X1 _5912_ (.A1(_1297_),
    .A2(net19),
    .ZN(_0047_));
 NOR2_X1 _5913_ (.A1(rst),
    .A2(net7),
    .ZN(_0046_));
 AND2_X1 _5914_ (.A1(_1297_),
    .A2(net33),
    .ZN(_0045_));
 NOR2_X1 _5915_ (.A1(rst),
    .A2(net52),
    .ZN(_0044_));
 AND2_X1 _5916_ (.A1(_1297_),
    .A2(net39),
    .ZN(_0043_));
 NOR2_X1 _5917_ (.A1(rst),
    .A2(net25),
    .ZN(_0042_));
 NOR2_X1 _5918_ (.A1(rst),
    .A2(net22),
    .ZN(_0041_));
 NOR2_X1 _5919_ (.A1(rst),
    .A2(net44),
    .ZN(_0040_));
 NOR2_X1 _5920_ (.A1(rst),
    .A2(net46),
    .ZN(_0039_));
 AND2_X1 _5921_ (.A1(_1297_),
    .A2(net31),
    .ZN(_0038_));
 AND2_X1 _5922_ (.A1(_1297_),
    .A2(net13),
    .ZN(_0037_));
 AND2_X1 _5923_ (.A1(_1297_),
    .A2(net41),
    .ZN(_0036_));
 AND2_X1 _5924_ (.A1(_1297_),
    .A2(net27),
    .ZN(_0035_));
 AND2_X1 _5925_ (.A1(_1297_),
    .A2(net15),
    .ZN(_0034_));
 AND2_X1 _5926_ (.A1(_1297_),
    .A2(net29),
    .ZN(_0033_));
 AND2_X1 _5927_ (.A1(_1297_),
    .A2(net35),
    .ZN(_0032_));
 DFF_X1 \iir1.t1[0]$_SDFF_PP0_  (.D(net36),
    .CK(clknet_3_7__leaf_clk),
    .Q(\iir1.t1[0] ),
    .QN(_3007_));
 DFF_X1 \iir1.t1[1]$_SDFF_PP0_  (.D(net30),
    .CK(clknet_3_7__leaf_clk),
    .Q(\iir1.t1[1] ),
    .QN(_3006_));
 DFF_X1 \iir1.t1[2]$_SDFF_PP0_  (.D(net16),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.t1[2] ),
    .QN(_3005_));
 DFF_X1 \iir1.t1[3]$_SDFF_PP0_  (.D(net28),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.t1[3] ),
    .QN(_3004_));
 DFF_X1 \iir1.t1[4]$_SDFF_PP0_  (.D(net42),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.t1[4] ),
    .QN(_3003_));
 DFF_X1 \iir1.x1[10]$_SDFF_PP0_  (.D(net14),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.x1[10] ),
    .QN(_3002_));
 DFF_X1 \iir1.x1[5]$_SDFF_PP0_  (.D(net32),
    .CK(clknet_3_4__leaf_clk),
    .Q(\iir1.x1[5] ),
    .QN(_3001_));
 DFF_X1 \iir1.x1[6]$_SDFF_PP0_  (.D(_0039_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\iir1.x1[6] ),
    .QN(_3000_));
 DFF_X1 \iir1.x1[7]$_SDFF_PP0_  (.D(_0040_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\iir1.x1[7] ),
    .QN(_2999_));
 DFF_X1 \iir1.x1[8]$_SDFF_PP0_  (.D(net23),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.x1[8] ),
    .QN(_2998_));
 DFF_X1 \iir1.x1[9]$_SDFF_PP0_  (.D(net26),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.x1[9] ),
    .QN(_2997_));
 DFF_X1 \iir1.x2[0]$_SDFF_PP0_  (.D(net40),
    .CK(clknet_3_6__leaf_clk),
    .Q(\iir1.x2[0] ),
    .QN(_2996_));
 DFF_X1 \iir1.x2[10]$_SDFF_PP0_  (.D(_0044_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.x2[10] ),
    .QN(_2995_));
 DFF_X1 \iir1.x2[1]$_SDFF_PP0_  (.D(net34),
    .CK(clknet_3_7__leaf_clk),
    .Q(\iir1.x2[1] ),
    .QN(_2994_));
 DFF_X1 \iir1.x2[2]$_SDFF_PP0_  (.D(net8),
    .CK(clknet_3_7__leaf_clk),
    .Q(\iir1.x2[2] ),
    .QN(_2993_));
 DFF_X1 \iir1.x2[3]$_SDFF_PP0_  (.D(net20),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.x2[3] ),
    .QN(_2992_));
 DFF_X1 \iir1.x2[4]$_SDFF_PP0_  (.D(net5),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.x2[4] ),
    .QN(_2991_));
 DFF_X1 \iir1.x2[5]$_SDFF_PP0_  (.D(net38),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.x2[5] ),
    .QN(_2990_));
 DFF_X1 \iir1.x2[6]$_SDFF_PP0_  (.D(net3),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.x2[6] ),
    .QN(_2989_));
 DFF_X1 \iir1.x2[7]$_SDFF_PP0_  (.D(net18),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.x2[7] ),
    .QN(_2988_));
 DFF_X1 \iir1.x2[8]$_SDFF_PP0_  (.D(net10),
    .CK(clknet_3_4__leaf_clk),
    .Q(\iir1.x2[8] ),
    .QN(_2987_));
 DFF_X1 \iir1.x2[9]$_SDFF_PP0_  (.D(net12),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.x2[9] ),
    .QN(_2986_));
 DFF_X1 \iir1.x[0]$_SDFF_PP0_  (.D(_0054_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\iir1.x[0] ),
    .QN(_2985_));
 DFF_X1 \iir1.x[10]$_SDFF_PP0_  (.D(_0055_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.x[10] ),
    .QN(_0010_));
 DFF_X1 \iir1.x[1]$_SDFF_PP0_  (.D(_0056_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\iir1.x[1] ),
    .QN(_2984_));
 DFF_X1 \iir1.x[2]$_SDFF_PP0_  (.D(_0057_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.x[2] ),
    .QN(_2983_));
 DFF_X1 \iir1.x[3]$_SDFF_PP0_  (.D(_0058_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\iir1.x[3] ),
    .QN(_2982_));
 DFF_X1 \iir1.x[4]$_SDFF_PP0_  (.D(_0059_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.x[4] ),
    .QN(_2981_));
 DFF_X1 \iir1.x[5]$_SDFF_PP0_  (.D(_0060_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\iir1.x[5] ),
    .QN(_2980_));
 DFF_X1 \iir1.x[6]$_SDFF_PP0_  (.D(_0061_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\iir1.x[6] ),
    .QN(_2979_));
 DFF_X1 \iir1.x[7]$_SDFF_PP0_  (.D(_0062_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\iir1.x[7] ),
    .QN(_2978_));
 DFF_X1 \iir1.x[8]$_SDFF_PP0_  (.D(_0063_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\iir1.x[8] ),
    .QN(_2977_));
 DFF_X1 \iir1.x[9]$_SDFF_PP0_  (.D(_0064_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\iir1.x[9] ),
    .QN(_2976_));
 DFF_X1 \iir1.y2[0]$_SDFF_PP0_  (.D(_0065_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\iir1.y2[0] ),
    .QN(_0015_));
 DFF_X1 \iir1.y2[10]$_SDFF_PP0_  (.D(net79),
    .CK(clknet_3_4__leaf_clk),
    .Q(\iir1.y2[10] ),
    .QN(_0004_));
 DFF_X1 \iir1.y2[1]$_SDFF_PP0_  (.D(_0067_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\iir1.y2[1] ),
    .QN(_0014_));
 DFF_X1 \iir1.y2[2]$_SDFF_PP0_  (.D(_0068_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\iir1.y2[2] ),
    .QN(_0013_));
 DFF_X1 \iir1.y2[3]$_SDFF_PP0_  (.D(_0069_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\iir1.y2[3] ),
    .QN(_0012_));
 DFF_X1 \iir1.y2[4]$_SDFF_PP0_  (.D(_0070_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\iir1.y2[4] ),
    .QN(_0011_));
 DFF_X1 \iir1.y2[5]$_SDFF_PP0_  (.D(_0071_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\iir1.y2[5] ),
    .QN(_0009_));
 DFF_X1 \iir1.y2[6]$_SDFF_PP0_  (.D(_0072_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\iir1.y2[6] ),
    .QN(_0003_));
 DFF_X1 \iir1.y2[7]$_SDFF_PP0_  (.D(_0073_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\iir1.y2[7] ),
    .QN(_0001_));
 DFF_X1 \iir1.y2[8]$_SDFF_PP0_  (.D(_0074_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\iir1.y2[8] ),
    .QN(_0008_));
 DFF_X1 \iir1.y2[9]$_SDFF_PP0_  (.D(net60),
    .CK(clknet_3_4__leaf_clk),
    .Q(\iir1.y2[9] ),
    .QN(_0030_));
 DFF_X1 \iir1.y[0]$_SDFF_PP0_  (.D(_0076_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\iir1.y[0] ),
    .QN(_2975_));
 DFF_X1 \iir1.y[10]$_SDFF_PP0_  (.D(_0077_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\iir1.y[10] ),
    .QN(_0006_));
 DFF_X1 \iir1.y[1]$_SDFF_PP0_  (.D(_0078_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\iir1.y[1] ),
    .QN(_2974_));
 DFF_X1 \iir1.y[2]$_SDFF_PP0_  (.D(_0079_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\iir1.y[2] ),
    .QN(_2973_));
 DFF_X1 \iir1.y[3]$_SDFF_PP0_  (.D(_0080_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\iir1.y[3] ),
    .QN(_2972_));
 DFF_X1 \iir1.y[4]$_SDFF_PP0_  (.D(_0081_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\iir1.y[4] ),
    .QN(_2971_));
 DFF_X1 \iir1.y[5]$_SDFF_PP0_  (.D(_0082_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\iir1.y[5] ),
    .QN(_0007_));
 DFF_X1 \iir1.y[6]$_SDFF_PP0_  (.D(_0083_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\iir1.y[6] ),
    .QN(_2970_));
 DFF_X1 \iir1.y[7]$_SDFF_PP0_  (.D(_0084_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\iir1.y[7] ),
    .QN(_2969_));
 DFF_X1 \iir1.y[8]$_SDFF_PP0_  (.D(_0085_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\iir1.y[8] ),
    .QN(_0005_));
 DFF_X1 \iir1.y[9]$_SDFF_PP0_  (.D(_0086_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\iir1.y[9] ),
    .QN(_0000_));
 DFF_X1 \iir2.x2[0]$_SDFF_PP0_  (.D(_0087_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\iir2.x2[0] ),
    .QN(_0024_));
 DFF_X1 \iir2.x2[10]$_SDFF_PP0_  (.D(_0088_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\iir2.x2[10] ),
    .QN(_0031_));
 DFF_X1 \iir2.x2[1]$_SDFF_PP0_  (.D(_0089_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\iir2.x2[1] ),
    .QN(_0023_));
 DFF_X1 \iir2.x2[2]$_SDFF_PP0_  (.D(_0090_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\iir2.x2[2] ),
    .QN(_0022_));
 DFF_X1 \iir2.x2[3]$_SDFF_PP0_  (.D(_0091_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\iir2.x2[3] ),
    .QN(_0021_));
 DFF_X1 \iir2.x2[4]$_SDFF_PP0_  (.D(_0092_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\iir2.x2[4] ),
    .QN(_0019_));
 DFF_X1 \iir2.x2[5]$_SDFF_PP0_  (.D(_0093_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\iir2.x2[5] ),
    .QN(_0017_));
 DFF_X1 \iir2.x2[6]$_SDFF_PP0_  (.D(_0094_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\iir2.x2[6] ),
    .QN(_0020_));
 DFF_X1 \iir2.x2[7]$_SDFF_PP0_  (.D(_0095_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\iir2.x2[7] ),
    .QN(_0018_));
 DFF_X1 \iir2.x2[8]$_SDFF_PP0_  (.D(_0096_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\iir2.x2[8] ),
    .QN(_0016_));
 DFF_X1 \iir2.x2[9]$_SDFF_PP0_  (.D(_0097_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\iir2.x2[9] ),
    .QN(_2968_));
 DFF_X1 \iir2.y2[0]$_SDFF_PP0_  (.D(_0098_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\iir2.y2[0] ),
    .QN(_0029_));
 DFF_X1 \iir2.y2[10]$_SDFF_PP0_  (.D(_0099_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\iir2.y2[10] ),
    .QN(_0002_));
 DFF_X1 \iir2.y2[1]$_SDFF_PP0_  (.D(net54),
    .CK(clknet_3_2__leaf_clk),
    .Q(\iir2.y2[1] ),
    .QN(_0027_));
 DFF_X1 \iir2.y2[2]$_SDFF_PP0_  (.D(net66),
    .CK(clknet_3_2__leaf_clk),
    .Q(\iir2.y2[2] ),
    .QN(_0025_));
 DFF_X1 \iir2.y2[3]$_SDFF_PP0_  (.D(net56),
    .CK(clknet_3_3__leaf_clk),
    .Q(\iir2.y2[3] ),
    .QN(_2967_));
 DFF_X1 \iir2.y2[4]$_SDFF_PP0_  (.D(_0103_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\iir2.y2[4] ),
    .QN(_2966_));
 DFF_X1 \iir2.y2[5]$_SDFF_PP0_  (.D(net58),
    .CK(clknet_3_6__leaf_clk),
    .Q(\iir2.y2[5] ),
    .QN(_0028_));
 DFF_X1 \iir2.y2[6]$_SDFF_PP0_  (.D(net81),
    .CK(clknet_3_6__leaf_clk),
    .Q(\iir2.y2[6] ),
    .QN(_0026_));
 DFF_X1 \iir2.y2[7]$_SDFF_PP0_  (.D(net68),
    .CK(clknet_3_3__leaf_clk),
    .Q(\iir2.y2[7] ),
    .QN(_2965_));
 DFF_X1 \iir2.y2[8]$_SDFF_PP0_  (.D(_0107_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\iir2.y2[8] ),
    .QN(_2964_));
 DFF_X1 \iir2.y2[9]$_SDFF_PP0_  (.D(_0108_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\iir2.y2[9] ),
    .QN(_2963_));
 DFF_X1 \z[0]$_SDFF_PP0_  (.D(_0109_),
    .CK(clknet_3_3__leaf_clk),
    .Q(z[0]),
    .QN(_2962_));
 DFF_X1 \z[10]$_SDFF_PP0_  (.D(_0110_),
    .CK(clknet_3_7__leaf_clk),
    .Q(z[10]),
    .QN(_2961_));
 DFF_X1 \z[1]$_SDFF_PP0_  (.D(_0111_),
    .CK(clknet_3_3__leaf_clk),
    .Q(z[1]),
    .QN(_2960_));
 DFF_X1 \z[2]$_SDFF_PP0_  (.D(_0112_),
    .CK(clknet_3_3__leaf_clk),
    .Q(z[2]),
    .QN(_2959_));
 DFF_X1 \z[3]$_SDFF_PP0_  (.D(_0113_),
    .CK(clknet_3_6__leaf_clk),
    .Q(z[3]),
    .QN(_2958_));
 DFF_X1 \z[4]$_SDFF_PP0_  (.D(_0114_),
    .CK(clknet_3_7__leaf_clk),
    .Q(z[4]),
    .QN(_2957_));
 DFF_X1 \z[5]$_SDFF_PP0_  (.D(_0115_),
    .CK(clknet_3_7__leaf_clk),
    .Q(z[5]),
    .QN(_2956_));
 DFF_X1 \z[6]$_SDFF_PP0_  (.D(_0116_),
    .CK(clknet_3_7__leaf_clk),
    .Q(z[6]),
    .QN(_2955_));
 DFF_X1 \z[7]$_SDFF_PP0_  (.D(_0117_),
    .CK(clknet_3_7__leaf_clk),
    .Q(z[7]),
    .QN(_2954_));
 DFF_X1 \z[8]$_SDFF_PP0_  (.D(_0118_),
    .CK(clknet_3_7__leaf_clk),
    .Q(z[8]),
    .QN(_2953_));
 DFF_X1 \z[9]$_SDFF_PP0_  (.D(_0119_),
    .CK(clknet_3_7__leaf_clk),
    .Q(z[9]),
    .QN(_2952_));
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_211 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_210 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_209 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_208 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_207 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_206 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_205 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_204 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_203 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_202 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_201 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_200 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_199 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_198 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_197 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_196 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_195 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_194 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_193 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_192 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_191 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_190 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_189 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_188 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_187 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_186 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_185 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_184 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_183 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_182 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_181 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_180 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_179 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_178 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_177 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_176 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_175 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_174 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_173 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_172 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_171 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_170 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_169 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_168 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_167 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_166 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_165 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_164 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_163 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_162 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_161 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_160 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_159 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_158 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_157 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_156 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_155 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_154 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_153 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_152 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_151 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_150 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_149 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_148 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_147 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_146 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_145 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_144 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_143 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_142 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_141 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_140 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_139 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_138 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_137 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_136 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_135 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_134 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_133 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_132 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_131 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_130 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_129 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_128 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_127 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_126 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_125 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_124 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_123 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_122 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_121 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_120 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_119 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_118 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_117 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_116 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_115 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_114 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_113 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_112 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_111 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_110 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_109 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_108 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_107 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_106 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_105 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_104 ();
 CLKBUF_X1 hold1 (.A(\iir1.x1[6] ),
    .Z(net1));
 CLKBUF_X1 hold2 (.A(_1233_),
    .Z(net2));
 CLKBUF_X1 hold3 (.A(_0050_),
    .Z(net3));
 CLKBUF_X1 hold4 (.A(net95),
    .Z(net4));
 CLKBUF_X1 hold5 (.A(_0048_),
    .Z(net5));
 CLKBUF_X1 hold6 (.A(\iir1.t1[2] ),
    .Z(net6));
 CLKBUF_X1 hold7 (.A(_1162_),
    .Z(net7));
 CLKBUF_X1 hold8 (.A(_0046_),
    .Z(net8));
 CLKBUF_X1 hold9 (.A(net96),
    .Z(net9));
 CLKBUF_X1 hold10 (.A(_0052_),
    .Z(net10));
 CLKBUF_X1 hold11 (.A(net97),
    .Z(net11));
 CLKBUF_X1 hold12 (.A(_0053_),
    .Z(net12));
 CLKBUF_X1 hold13 (.A(net98),
    .Z(net13));
 CLKBUF_X1 hold14 (.A(_0037_),
    .Z(net14));
 CLKBUF_X1 hold15 (.A(net99),
    .Z(net15));
 CLKBUF_X1 hold16 (.A(_0034_),
    .Z(net16));
 CLKBUF_X1 hold17 (.A(net100),
    .Z(net17));
 CLKBUF_X1 hold18 (.A(_0051_),
    .Z(net18));
 CLKBUF_X1 hold19 (.A(net101),
    .Z(net19));
 CLKBUF_X1 hold20 (.A(_0047_),
    .Z(net20));
 CLKBUF_X1 hold21 (.A(\iir1.x[8] ),
    .Z(net21));
 CLKBUF_X1 hold22 (.A(_1022_),
    .Z(net22));
 CLKBUF_X1 hold23 (.A(_0041_),
    .Z(net23));
 CLKBUF_X1 hold24 (.A(\iir1.x[9] ),
    .Z(net24));
 CLKBUF_X1 hold25 (.A(_1230_),
    .Z(net25));
 CLKBUF_X1 hold26 (.A(_0042_),
    .Z(net26));
 CLKBUF_X1 hold27 (.A(net102),
    .Z(net27));
 CLKBUF_X1 hold28 (.A(_0035_),
    .Z(net28));
 CLKBUF_X1 hold29 (.A(net103),
    .Z(net29));
 CLKBUF_X1 hold30 (.A(_0033_),
    .Z(net30));
 CLKBUF_X1 hold31 (.A(net107),
    .Z(net31));
 CLKBUF_X1 hold32 (.A(_0038_),
    .Z(net32));
 CLKBUF_X1 hold33 (.A(net104),
    .Z(net33));
 CLKBUF_X1 hold34 (.A(_0045_),
    .Z(net34));
 CLKBUF_X1 hold35 (.A(net106),
    .Z(net35));
 CLKBUF_X1 hold36 (.A(_0032_),
    .Z(net36));
 CLKBUF_X1 hold37 (.A(net105),
    .Z(net37));
 CLKBUF_X1 hold38 (.A(_0049_),
    .Z(net38));
 CLKBUF_X1 hold39 (.A(net111),
    .Z(net39));
 CLKBUF_X1 hold40 (.A(_0043_),
    .Z(net40));
 CLKBUF_X1 hold41 (.A(net109),
    .Z(net41));
 CLKBUF_X1 hold42 (.A(_0036_),
    .Z(net42));
 CLKBUF_X1 hold43 (.A(net118),
    .Z(net43));
 CLKBUF_X1 hold44 (.A(_0947_),
    .Z(net44));
 CLKBUF_X1 hold45 (.A(\iir1.x[6] ),
    .Z(net45));
 CLKBUF_X1 hold46 (.A(_0917_),
    .Z(net46));
 CLKBUF_X1 hold47 (.A(net125),
    .Z(net47));
 CLKBUF_X1 hold48 (.A(_2385_),
    .Z(net48));
 CLKBUF_X1 hold49 (.A(z[0]),
    .Z(net49));
 CLKBUF_X1 hold50 (.A(_2849_),
    .Z(net50));
 CLKBUF_X1 hold51 (.A(\iir1.x1[10] ),
    .Z(net51));
 CLKBUF_X1 hold52 (.A(_1592_),
    .Z(net52));
 CLKBUF_X1 hold53 (.A(net122),
    .Z(net53));
 CLKBUF_X1 hold54 (.A(_0100_),
    .Z(net54));
 CLKBUF_X1 hold55 (.A(z[3]),
    .Z(net55));
 CLKBUF_X1 hold56 (.A(_0102_),
    .Z(net56));
 CLKBUF_X1 hold57 (.A(z[5]),
    .Z(net57));
 CLKBUF_X1 hold58 (.A(_0104_),
    .Z(net58));
 CLKBUF_X1 hold59 (.A(net126),
    .Z(net59));
 CLKBUF_X1 hold60 (.A(_0075_),
    .Z(net60));
 CLKBUF_X1 hold61 (.A(\iir1.y2[6] ),
    .Z(net61));
 CLKBUF_X1 hold62 (.A(_2430_),
    .Z(net62));
 CLKBUF_X1 hold63 (.A(z[9]),
    .Z(net63));
 CLKBUF_X1 hold64 (.A(_2753_),
    .Z(net64));
 CLKBUF_X1 hold65 (.A(z[2]),
    .Z(net65));
 CLKBUF_X1 hold66 (.A(_0101_),
    .Z(net66));
 CLKBUF_X1 hold67 (.A(z[7]),
    .Z(net67));
 CLKBUF_X1 hold68 (.A(_0106_),
    .Z(net68));
 CLKBUF_X1 hold69 (.A(net108),
    .Z(net69));
 CLKBUF_X1 hold70 (.A(\iir1.y2[8] ),
    .Z(net70));
 CLKBUF_X1 hold71 (.A(_2491_),
    .Z(net71));
 CLKBUF_X1 hold72 (.A(\iir1.y2[3] ),
    .Z(net72));
 CLKBUF_X1 hold73 (.A(_0906_),
    .Z(net73));
 CLKBUF_X1 hold74 (.A(net112),
    .Z(net74));
 CLKBUF_X1 hold75 (.A(net110),
    .Z(net75));
 CLKBUF_X1 hold76 (.A(\iir1.y2[2] ),
    .Z(net76));
 CLKBUF_X1 hold77 (.A(_1506_),
    .Z(net77));
 CLKBUF_X1 hold78 (.A(\iir1.y[10] ),
    .Z(net78));
 CLKBUF_X1 hold79 (.A(_0066_),
    .Z(net79));
 CLKBUF_X1 hold80 (.A(z[6]),
    .Z(net80));
 CLKBUF_X1 hold81 (.A(_0105_),
    .Z(net81));
 CLKBUF_X1 hold82 (.A(net113),
    .Z(net82));
 CLKBUF_X1 hold83 (.A(net114),
    .Z(net83));
 CLKBUF_X1 hold84 (.A(net115),
    .Z(net84));
 CLKBUF_X1 hold85 (.A(net117),
    .Z(net85));
 CLKBUF_X1 hold86 (.A(net119),
    .Z(net86));
 CLKBUF_X1 hold87 (.A(net116),
    .Z(net87));
 CLKBUF_X1 hold88 (.A(net120),
    .Z(net88));
 CLKBUF_X1 hold89 (.A(net121),
    .Z(net89));
 CLKBUF_X1 hold90 (.A(net123),
    .Z(net90));
 CLKBUF_X1 hold91 (.A(net124),
    .Z(net91));
 CLKBUF_X1 hold92 (.A(\iir1.y[6] ),
    .Z(net92));
 CLKBUF_X1 hold93 (.A(\iir1.y[1] ),
    .Z(net93));
 CLKBUF_X1 hold94 (.A(\iir1.y[7] ),
    .Z(net94));
 CLKBUF_X1 hold95 (.A(\iir1.t1[4] ),
    .Z(net95));
 CLKBUF_X1 hold96 (.A(\iir1.x1[8] ),
    .Z(net96));
 CLKBUF_X1 hold97 (.A(\iir1.x1[9] ),
    .Z(net97));
 CLKBUF_X1 hold98 (.A(\iir1.x[10] ),
    .Z(net98));
 CLKBUF_X1 hold99 (.A(\iir1.x[2] ),
    .Z(net99));
 CLKBUF_X1 hold100 (.A(\iir1.x1[7] ),
    .Z(net100));
 CLKBUF_X1 hold101 (.A(\iir1.t1[3] ),
    .Z(net101));
 CLKBUF_X1 hold102 (.A(\iir1.x[3] ),
    .Z(net102));
 CLKBUF_X1 hold103 (.A(\iir1.x[1] ),
    .Z(net103));
 CLKBUF_X1 hold104 (.A(\iir1.t1[1] ),
    .Z(net104));
 CLKBUF_X1 hold105 (.A(\iir1.x1[5] ),
    .Z(net105));
 CLKBUF_X1 hold106 (.A(\iir1.x[0] ),
    .Z(net106));
 CLKBUF_X1 hold107 (.A(\iir1.x[5] ),
    .Z(net107));
 BUF_X8 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 BUF_X8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk));
 BUF_X8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk));
 BUF_X8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk));
 BUF_X8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk));
 BUF_X8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk));
 BUF_X8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk));
 BUF_X8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk));
 BUF_X8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk));
 BUF_X8 clkload0 (.A(clknet_3_0__leaf_clk));
 INV_X8 clkload1 (.A(clknet_3_1__leaf_clk));
 BUF_X4 clkload2 (.A(clknet_3_2__leaf_clk));
 BUF_X8 clkload3 (.A(clknet_3_3__leaf_clk));
 BUF_X4 clkload4 (.A(clknet_3_4__leaf_clk));
 BUF_X8 clkload5 (.A(clknet_3_6__leaf_clk));
 BUF_X4 clkload6 (.A(clknet_3_7__leaf_clk));
 CLKBUF_X1 hold108 (.A(z[4]),
    .Z(net108));
 CLKBUF_X1 hold109 (.A(\iir1.x[4] ),
    .Z(net109));
 CLKBUF_X1 hold110 (.A(z[10]),
    .Z(net110));
 CLKBUF_X1 hold111 (.A(\iir1.t1[0] ),
    .Z(net111));
 CLKBUF_X1 hold112 (.A(z[8]),
    .Z(net112));
 CLKBUF_X1 hold113 (.A(\iir1.y2[4] ),
    .Z(net113));
 CLKBUF_X1 hold114 (.A(\iir1.y[8] ),
    .Z(net114));
 CLKBUF_X1 hold115 (.A(\iir1.y2[1] ),
    .Z(net115));
 CLKBUF_X1 hold116 (.A(\iir1.y2[9] ),
    .Z(net116));
 CLKBUF_X1 hold117 (.A(\iir1.y2[7] ),
    .Z(net117));
 CLKBUF_X1 hold118 (.A(\iir1.x[7] ),
    .Z(net118));
 CLKBUF_X1 hold119 (.A(\iir1.y[5] ),
    .Z(net119));
 CLKBUF_X1 hold120 (.A(\iir1.y2[5] ),
    .Z(net120));
 CLKBUF_X1 hold121 (.A(\iir1.y[4] ),
    .Z(net121));
 CLKBUF_X1 hold122 (.A(z[1]),
    .Z(net122));
 CLKBUF_X1 hold123 (.A(\iir1.y[2] ),
    .Z(net123));
 CLKBUF_X1 hold124 (.A(\iir1.y[3] ),
    .Z(net124));
 CLKBUF_X1 hold125 (.A(\iir1.y2[0] ),
    .Z(net125));
 CLKBUF_X1 hold126 (.A(\iir1.y[9] ),
    .Z(net126));
 FILLCELL_X32 FILLER_0_0_1 ();
 FILLCELL_X8 FILLER_0_0_33 ();
 FILLCELL_X8 FILLER_0_0_51 ();
 FILLCELL_X4 FILLER_0_0_77 ();
 FILLCELL_X2 FILLER_0_0_81 ();
 FILLCELL_X2 FILLER_0_0_90 ();
 FILLCELL_X2 FILLER_0_0_98 ();
 FILLCELL_X1 FILLER_0_0_100 ();
 FILLCELL_X8 FILLER_0_0_114 ();
 FILLCELL_X2 FILLER_0_0_122 ();
 FILLCELL_X1 FILLER_0_0_124 ();
 FILLCELL_X2 FILLER_0_0_128 ();
 FILLCELL_X1 FILLER_0_0_130 ();
 FILLCELL_X1 FILLER_0_0_135 ();
 FILLCELL_X1 FILLER_0_0_142 ();
 FILLCELL_X8 FILLER_0_0_146 ();
 FILLCELL_X8 FILLER_0_0_159 ();
 FILLCELL_X1 FILLER_0_0_167 ();
 FILLCELL_X2 FILLER_0_0_172 ();
 FILLCELL_X1 FILLER_0_0_174 ();
 FILLCELL_X4 FILLER_0_0_183 ();
 FILLCELL_X2 FILLER_0_0_187 ();
 FILLCELL_X1 FILLER_0_0_189 ();
 FILLCELL_X1 FILLER_0_0_205 ();
 FILLCELL_X2 FILLER_0_0_215 ();
 FILLCELL_X1 FILLER_0_0_217 ();
 FILLCELL_X16 FILLER_0_0_222 ();
 FILLCELL_X8 FILLER_0_0_238 ();
 FILLCELL_X1 FILLER_0_0_246 ();
 FILLCELL_X2 FILLER_0_0_256 ();
 FILLCELL_X1 FILLER_0_0_258 ();
 FILLCELL_X2 FILLER_0_0_261 ();
 FILLCELL_X8 FILLER_0_0_268 ();
 FILLCELL_X2 FILLER_0_0_276 ();
 FILLCELL_X1 FILLER_0_0_278 ();
 FILLCELL_X4 FILLER_0_0_289 ();
 FILLCELL_X4 FILLER_0_0_297 ();
 FILLCELL_X2 FILLER_0_0_315 ();
 FILLCELL_X1 FILLER_0_0_317 ();
 FILLCELL_X4 FILLER_0_0_324 ();
 FILLCELL_X2 FILLER_0_0_342 ();
 FILLCELL_X2 FILLER_0_0_348 ();
 FILLCELL_X1 FILLER_0_0_350 ();
 FILLCELL_X1 FILLER_0_0_355 ();
 FILLCELL_X8 FILLER_0_0_362 ();
 FILLCELL_X2 FILLER_0_0_370 ();
 FILLCELL_X1 FILLER_0_0_372 ();
 FILLCELL_X8 FILLER_0_0_377 ();
 FILLCELL_X2 FILLER_0_0_385 ();
 FILLCELL_X1 FILLER_0_0_387 ();
 FILLCELL_X32 FILLER_0_1_1 ();
 FILLCELL_X4 FILLER_0_1_33 ();
 FILLCELL_X2 FILLER_0_1_37 ();
 FILLCELL_X1 FILLER_0_1_39 ();
 FILLCELL_X4 FILLER_0_1_54 ();
 FILLCELL_X1 FILLER_0_1_58 ();
 FILLCELL_X1 FILLER_0_1_65 ();
 FILLCELL_X1 FILLER_0_1_70 ();
 FILLCELL_X1 FILLER_0_1_77 ();
 FILLCELL_X2 FILLER_0_1_84 ();
 FILLCELL_X2 FILLER_0_1_96 ();
 FILLCELL_X1 FILLER_0_1_98 ();
 FILLCELL_X2 FILLER_0_1_102 ();
 FILLCELL_X1 FILLER_0_1_104 ();
 FILLCELL_X1 FILLER_0_1_127 ();
 FILLCELL_X1 FILLER_0_1_140 ();
 FILLCELL_X1 FILLER_0_1_144 ();
 FILLCELL_X8 FILLER_0_1_162 ();
 FILLCELL_X2 FILLER_0_1_170 ();
 FILLCELL_X1 FILLER_0_1_190 ();
 FILLCELL_X2 FILLER_0_1_208 ();
 FILLCELL_X2 FILLER_0_1_216 ();
 FILLCELL_X1 FILLER_0_1_224 ();
 FILLCELL_X8 FILLER_0_1_228 ();
 FILLCELL_X4 FILLER_0_1_242 ();
 FILLCELL_X2 FILLER_0_1_250 ();
 FILLCELL_X1 FILLER_0_1_252 ();
 FILLCELL_X2 FILLER_0_1_277 ();
 FILLCELL_X1 FILLER_0_1_313 ();
 FILLCELL_X2 FILLER_0_1_318 ();
 FILLCELL_X1 FILLER_0_1_330 ();
 FILLCELL_X1 FILLER_0_1_335 ();
 FILLCELL_X1 FILLER_0_1_345 ();
 FILLCELL_X1 FILLER_0_1_355 ();
 FILLCELL_X8 FILLER_0_1_357 ();
 FILLCELL_X4 FILLER_0_1_365 ();
 FILLCELL_X1 FILLER_0_1_369 ();
 FILLCELL_X1 FILLER_0_1_387 ();
 FILLCELL_X32 FILLER_0_2_1 ();
 FILLCELL_X1 FILLER_0_2_33 ();
 FILLCELL_X4 FILLER_0_2_64 ();
 FILLCELL_X1 FILLER_0_2_78 ();
 FILLCELL_X1 FILLER_0_2_88 ();
 FILLCELL_X1 FILLER_0_2_90 ();
 FILLCELL_X1 FILLER_0_2_97 ();
 FILLCELL_X1 FILLER_0_2_102 ();
 FILLCELL_X1 FILLER_0_2_109 ();
 FILLCELL_X1 FILLER_0_2_133 ();
 FILLCELL_X2 FILLER_0_2_149 ();
 FILLCELL_X8 FILLER_0_2_176 ();
 FILLCELL_X1 FILLER_0_2_184 ();
 FILLCELL_X2 FILLER_0_2_194 ();
 FILLCELL_X2 FILLER_0_2_215 ();
 FILLCELL_X4 FILLER_0_2_227 ();
 FILLCELL_X1 FILLER_0_2_231 ();
 FILLCELL_X4 FILLER_0_2_249 ();
 FILLCELL_X1 FILLER_0_2_253 ();
 FILLCELL_X1 FILLER_0_2_266 ();
 FILLCELL_X4 FILLER_0_2_268 ();
 FILLCELL_X1 FILLER_0_2_285 ();
 FILLCELL_X8 FILLER_0_2_290 ();
 FILLCELL_X1 FILLER_0_2_298 ();
 FILLCELL_X2 FILLER_0_2_305 ();
 FILLCELL_X2 FILLER_0_2_313 ();
 FILLCELL_X1 FILLER_0_2_315 ();
 FILLCELL_X1 FILLER_0_2_362 ();
 FILLCELL_X16 FILLER_0_2_369 ();
 FILLCELL_X2 FILLER_0_2_385 ();
 FILLCELL_X1 FILLER_0_2_387 ();
 FILLCELL_X16 FILLER_0_3_1 ();
 FILLCELL_X8 FILLER_0_3_17 ();
 FILLCELL_X4 FILLER_0_3_25 ();
 FILLCELL_X2 FILLER_0_3_29 ();
 FILLCELL_X1 FILLER_0_3_31 ();
 FILLCELL_X2 FILLER_0_3_41 ();
 FILLCELL_X1 FILLER_0_3_54 ();
 FILLCELL_X4 FILLER_0_3_65 ();
 FILLCELL_X1 FILLER_0_3_93 ();
 FILLCELL_X1 FILLER_0_3_104 ();
 FILLCELL_X1 FILLER_0_3_109 ();
 FILLCELL_X4 FILLER_0_3_119 ();
 FILLCELL_X1 FILLER_0_3_123 ();
 FILLCELL_X4 FILLER_0_3_164 ();
 FILLCELL_X2 FILLER_0_3_168 ();
 FILLCELL_X2 FILLER_0_3_176 ();
 FILLCELL_X4 FILLER_0_3_179 ();
 FILLCELL_X1 FILLER_0_3_183 ();
 FILLCELL_X2 FILLER_0_3_210 ();
 FILLCELL_X1 FILLER_0_3_231 ();
 FILLCELL_X1 FILLER_0_3_236 ();
 FILLCELL_X1 FILLER_0_3_254 ();
 FILLCELL_X1 FILLER_0_3_265 ();
 FILLCELL_X2 FILLER_0_3_275 ();
 FILLCELL_X1 FILLER_0_3_286 ();
 FILLCELL_X2 FILLER_0_3_303 ();
 FILLCELL_X1 FILLER_0_3_305 ();
 FILLCELL_X2 FILLER_0_3_319 ();
 FILLCELL_X1 FILLER_0_3_321 ();
 FILLCELL_X1 FILLER_0_3_343 ();
 FILLCELL_X4 FILLER_0_3_350 ();
 FILLCELL_X2 FILLER_0_3_354 ();
 FILLCELL_X2 FILLER_0_3_357 ();
 FILLCELL_X2 FILLER_0_3_379 ();
 FILLCELL_X4 FILLER_0_3_384 ();
 FILLCELL_X16 FILLER_0_4_1 ();
 FILLCELL_X8 FILLER_0_4_17 ();
 FILLCELL_X1 FILLER_0_4_50 ();
 FILLCELL_X2 FILLER_0_4_55 ();
 FILLCELL_X4 FILLER_0_4_60 ();
 FILLCELL_X2 FILLER_0_4_64 ();
 FILLCELL_X1 FILLER_0_4_66 ();
 FILLCELL_X1 FILLER_0_4_76 ();
 FILLCELL_X2 FILLER_0_4_105 ();
 FILLCELL_X1 FILLER_0_4_113 ();
 FILLCELL_X8 FILLER_0_4_118 ();
 FILLCELL_X2 FILLER_0_4_126 ();
 FILLCELL_X1 FILLER_0_4_128 ();
 FILLCELL_X8 FILLER_0_4_138 ();
 FILLCELL_X2 FILLER_0_4_146 ();
 FILLCELL_X1 FILLER_0_4_148 ();
 FILLCELL_X1 FILLER_0_4_173 ();
 FILLCELL_X1 FILLER_0_4_187 ();
 FILLCELL_X1 FILLER_0_4_213 ();
 FILLCELL_X8 FILLER_0_4_237 ();
 FILLCELL_X4 FILLER_0_4_245 ();
 FILLCELL_X1 FILLER_0_4_249 ();
 FILLCELL_X4 FILLER_0_4_259 ();
 FILLCELL_X1 FILLER_0_4_268 ();
 FILLCELL_X1 FILLER_0_4_272 ();
 FILLCELL_X1 FILLER_0_4_278 ();
 FILLCELL_X1 FILLER_0_4_285 ();
 FILLCELL_X1 FILLER_0_4_288 ();
 FILLCELL_X1 FILLER_0_4_295 ();
 FILLCELL_X1 FILLER_0_4_299 ();
 FILLCELL_X2 FILLER_0_4_306 ();
 FILLCELL_X4 FILLER_0_4_313 ();
 FILLCELL_X2 FILLER_0_4_325 ();
 FILLCELL_X1 FILLER_0_4_327 ();
 FILLCELL_X1 FILLER_0_4_331 ();
 FILLCELL_X1 FILLER_0_4_339 ();
 FILLCELL_X8 FILLER_0_4_354 ();
 FILLCELL_X2 FILLER_0_4_369 ();
 FILLCELL_X8 FILLER_0_5_1 ();
 FILLCELL_X4 FILLER_0_5_9 ();
 FILLCELL_X2 FILLER_0_5_13 ();
 FILLCELL_X1 FILLER_0_5_15 ();
 FILLCELL_X2 FILLER_0_5_33 ();
 FILLCELL_X1 FILLER_0_5_38 ();
 FILLCELL_X2 FILLER_0_5_62 ();
 FILLCELL_X2 FILLER_0_5_73 ();
 FILLCELL_X4 FILLER_0_5_85 ();
 FILLCELL_X1 FILLER_0_5_92 ();
 FILLCELL_X16 FILLER_0_5_109 ();
 FILLCELL_X2 FILLER_0_5_125 ();
 FILLCELL_X1 FILLER_0_5_145 ();
 FILLCELL_X1 FILLER_0_5_156 ();
 FILLCELL_X1 FILLER_0_5_161 ();
 FILLCELL_X4 FILLER_0_5_167 ();
 FILLCELL_X1 FILLER_0_5_171 ();
 FILLCELL_X2 FILLER_0_5_179 ();
 FILLCELL_X2 FILLER_0_5_191 ();
 FILLCELL_X8 FILLER_0_5_195 ();
 FILLCELL_X1 FILLER_0_5_203 ();
 FILLCELL_X8 FILLER_0_5_237 ();
 FILLCELL_X4 FILLER_0_5_245 ();
 FILLCELL_X2 FILLER_0_5_288 ();
 FILLCELL_X1 FILLER_0_5_290 ();
 FILLCELL_X1 FILLER_0_5_294 ();
 FILLCELL_X1 FILLER_0_5_297 ();
 FILLCELL_X2 FILLER_0_5_308 ();
 FILLCELL_X1 FILLER_0_5_321 ();
 FILLCELL_X1 FILLER_0_5_339 ();
 FILLCELL_X1 FILLER_0_5_349 ();
 FILLCELL_X1 FILLER_0_5_377 ();
 FILLCELL_X8 FILLER_0_5_380 ();
 FILLCELL_X16 FILLER_0_6_1 ();
 FILLCELL_X2 FILLER_0_6_17 ();
 FILLCELL_X1 FILLER_0_6_38 ();
 FILLCELL_X1 FILLER_0_6_43 ();
 FILLCELL_X1 FILLER_0_6_48 ();
 FILLCELL_X1 FILLER_0_6_60 ();
 FILLCELL_X2 FILLER_0_6_67 ();
 FILLCELL_X1 FILLER_0_6_90 ();
 FILLCELL_X4 FILLER_0_6_101 ();
 FILLCELL_X1 FILLER_0_6_105 ();
 FILLCELL_X8 FILLER_0_6_108 ();
 FILLCELL_X2 FILLER_0_6_116 ();
 FILLCELL_X1 FILLER_0_6_146 ();
 FILLCELL_X2 FILLER_0_6_150 ();
 FILLCELL_X1 FILLER_0_6_161 ();
 FILLCELL_X1 FILLER_0_6_174 ();
 FILLCELL_X4 FILLER_0_6_179 ();
 FILLCELL_X1 FILLER_0_6_183 ();
 FILLCELL_X4 FILLER_0_6_204 ();
 FILLCELL_X2 FILLER_0_6_208 ();
 FILLCELL_X1 FILLER_0_6_210 ();
 FILLCELL_X8 FILLER_0_6_222 ();
 FILLCELL_X1 FILLER_0_6_230 ();
 FILLCELL_X1 FILLER_0_6_244 ();
 FILLCELL_X1 FILLER_0_6_254 ();
 FILLCELL_X1 FILLER_0_6_257 ();
 FILLCELL_X1 FILLER_0_6_272 ();
 FILLCELL_X2 FILLER_0_6_277 ();
 FILLCELL_X1 FILLER_0_6_279 ();
 FILLCELL_X2 FILLER_0_6_313 ();
 FILLCELL_X2 FILLER_0_6_324 ();
 FILLCELL_X1 FILLER_0_6_371 ();
 FILLCELL_X8 FILLER_0_6_380 ();
 FILLCELL_X8 FILLER_0_7_1 ();
 FILLCELL_X1 FILLER_0_7_9 ();
 FILLCELL_X8 FILLER_0_7_14 ();
 FILLCELL_X2 FILLER_0_7_22 ();
 FILLCELL_X4 FILLER_0_7_57 ();
 FILLCELL_X2 FILLER_0_7_61 ();
 FILLCELL_X4 FILLER_0_7_67 ();
 FILLCELL_X4 FILLER_0_7_77 ();
 FILLCELL_X4 FILLER_0_7_87 ();
 FILLCELL_X1 FILLER_0_7_97 ();
 FILLCELL_X1 FILLER_0_7_101 ();
 FILLCELL_X1 FILLER_0_7_105 ();
 FILLCELL_X2 FILLER_0_7_109 ();
 FILLCELL_X1 FILLER_0_7_140 ();
 FILLCELL_X2 FILLER_0_7_150 ();
 FILLCELL_X1 FILLER_0_7_161 ();
 FILLCELL_X1 FILLER_0_7_177 ();
 FILLCELL_X4 FILLER_0_7_179 ();
 FILLCELL_X1 FILLER_0_7_189 ();
 FILLCELL_X2 FILLER_0_7_216 ();
 FILLCELL_X16 FILLER_0_7_222 ();
 FILLCELL_X2 FILLER_0_7_247 ();
 FILLCELL_X2 FILLER_0_7_251 ();
 FILLCELL_X1 FILLER_0_7_253 ();
 FILLCELL_X2 FILLER_0_7_286 ();
 FILLCELL_X1 FILLER_0_7_291 ();
 FILLCELL_X1 FILLER_0_7_314 ();
 FILLCELL_X2 FILLER_0_7_318 ();
 FILLCELL_X1 FILLER_0_7_323 ();
 FILLCELL_X2 FILLER_0_7_327 ();
 FILLCELL_X4 FILLER_0_7_332 ();
 FILLCELL_X2 FILLER_0_7_336 ();
 FILLCELL_X1 FILLER_0_7_338 ();
 FILLCELL_X1 FILLER_0_7_365 ();
 FILLCELL_X4 FILLER_0_7_384 ();
 FILLCELL_X16 FILLER_0_8_1 ();
 FILLCELL_X8 FILLER_0_8_17 ();
 FILLCELL_X2 FILLER_0_8_25 ();
 FILLCELL_X1 FILLER_0_8_27 ();
 FILLCELL_X1 FILLER_0_8_52 ();
 FILLCELL_X1 FILLER_0_8_62 ();
 FILLCELL_X16 FILLER_0_8_69 ();
 FILLCELL_X4 FILLER_0_8_85 ();
 FILLCELL_X2 FILLER_0_8_90 ();
 FILLCELL_X1 FILLER_0_8_92 ();
 FILLCELL_X1 FILLER_0_8_121 ();
 FILLCELL_X2 FILLER_0_8_126 ();
 FILLCELL_X1 FILLER_0_8_128 ();
 FILLCELL_X4 FILLER_0_8_139 ();
 FILLCELL_X1 FILLER_0_8_143 ();
 FILLCELL_X2 FILLER_0_8_154 ();
 FILLCELL_X1 FILLER_0_8_156 ();
 FILLCELL_X1 FILLER_0_8_180 ();
 FILLCELL_X4 FILLER_0_8_184 ();
 FILLCELL_X4 FILLER_0_8_191 ();
 FILLCELL_X1 FILLER_0_8_195 ();
 FILLCELL_X2 FILLER_0_8_212 ();
 FILLCELL_X1 FILLER_0_8_214 ();
 FILLCELL_X16 FILLER_0_8_229 ();
 FILLCELL_X1 FILLER_0_8_261 ();
 FILLCELL_X1 FILLER_0_8_266 ();
 FILLCELL_X2 FILLER_0_8_294 ();
 FILLCELL_X1 FILLER_0_8_307 ();
 FILLCELL_X1 FILLER_0_8_325 ();
 FILLCELL_X2 FILLER_0_8_358 ();
 FILLCELL_X2 FILLER_0_8_386 ();
 FILLCELL_X4 FILLER_0_9_1 ();
 FILLCELL_X2 FILLER_0_9_5 ();
 FILLCELL_X1 FILLER_0_9_7 ();
 FILLCELL_X4 FILLER_0_9_48 ();
 FILLCELL_X1 FILLER_0_9_52 ();
 FILLCELL_X1 FILLER_0_9_70 ();
 FILLCELL_X1 FILLER_0_9_88 ();
 FILLCELL_X1 FILLER_0_9_95 ();
 FILLCELL_X1 FILLER_0_9_99 ();
 FILLCELL_X4 FILLER_0_9_119 ();
 FILLCELL_X2 FILLER_0_9_123 ();
 FILLCELL_X1 FILLER_0_9_125 ();
 FILLCELL_X2 FILLER_0_9_135 ();
 FILLCELL_X2 FILLER_0_9_161 ();
 FILLCELL_X2 FILLER_0_9_173 ();
 FILLCELL_X2 FILLER_0_9_185 ();
 FILLCELL_X1 FILLER_0_9_187 ();
 FILLCELL_X2 FILLER_0_9_228 ();
 FILLCELL_X8 FILLER_0_9_236 ();
 FILLCELL_X1 FILLER_0_9_244 ();
 FILLCELL_X2 FILLER_0_9_274 ();
 FILLCELL_X2 FILLER_0_9_279 ();
 FILLCELL_X1 FILLER_0_9_281 ();
 FILLCELL_X4 FILLER_0_9_288 ();
 FILLCELL_X2 FILLER_0_9_292 ();
 FILLCELL_X1 FILLER_0_9_307 ();
 FILLCELL_X1 FILLER_0_9_325 ();
 FILLCELL_X1 FILLER_0_9_329 ();
 FILLCELL_X2 FILLER_0_9_334 ();
 FILLCELL_X2 FILLER_0_9_366 ();
 FILLCELL_X1 FILLER_0_9_368 ();
 FILLCELL_X1 FILLER_0_9_387 ();
 FILLCELL_X4 FILLER_0_10_1 ();
 FILLCELL_X2 FILLER_0_10_5 ();
 FILLCELL_X1 FILLER_0_10_7 ();
 FILLCELL_X8 FILLER_0_10_29 ();
 FILLCELL_X2 FILLER_0_10_54 ();
 FILLCELL_X8 FILLER_0_10_60 ();
 FILLCELL_X4 FILLER_0_10_68 ();
 FILLCELL_X1 FILLER_0_10_113 ();
 FILLCELL_X1 FILLER_0_10_120 ();
 FILLCELL_X1 FILLER_0_10_131 ();
 FILLCELL_X4 FILLER_0_10_141 ();
 FILLCELL_X1 FILLER_0_10_145 ();
 FILLCELL_X2 FILLER_0_10_166 ();
 FILLCELL_X1 FILLER_0_10_185 ();
 FILLCELL_X1 FILLER_0_10_192 ();
 FILLCELL_X1 FILLER_0_10_208 ();
 FILLCELL_X8 FILLER_0_10_213 ();
 FILLCELL_X2 FILLER_0_10_241 ();
 FILLCELL_X1 FILLER_0_10_259 ();
 FILLCELL_X2 FILLER_0_10_264 ();
 FILLCELL_X1 FILLER_0_10_266 ();
 FILLCELL_X1 FILLER_0_10_280 ();
 FILLCELL_X1 FILLER_0_10_291 ();
 FILLCELL_X1 FILLER_0_10_298 ();
 FILLCELL_X1 FILLER_0_10_305 ();
 FILLCELL_X1 FILLER_0_10_309 ();
 FILLCELL_X2 FILLER_0_10_313 ();
 FILLCELL_X1 FILLER_0_10_331 ();
 FILLCELL_X4 FILLER_0_10_352 ();
 FILLCELL_X1 FILLER_0_10_356 ();
 FILLCELL_X4 FILLER_0_10_383 ();
 FILLCELL_X1 FILLER_0_10_387 ();
 FILLCELL_X4 FILLER_0_11_1 ();
 FILLCELL_X1 FILLER_0_11_29 ();
 FILLCELL_X2 FILLER_0_11_34 ();
 FILLCELL_X2 FILLER_0_11_47 ();
 FILLCELL_X4 FILLER_0_11_80 ();
 FILLCELL_X1 FILLER_0_11_84 ();
 FILLCELL_X1 FILLER_0_11_93 ();
 FILLCELL_X2 FILLER_0_11_100 ();
 FILLCELL_X4 FILLER_0_11_110 ();
 FILLCELL_X1 FILLER_0_11_114 ();
 FILLCELL_X1 FILLER_0_11_122 ();
 FILLCELL_X4 FILLER_0_11_132 ();
 FILLCELL_X4 FILLER_0_11_139 ();
 FILLCELL_X1 FILLER_0_11_143 ();
 FILLCELL_X4 FILLER_0_11_154 ();
 FILLCELL_X2 FILLER_0_11_158 ();
 FILLCELL_X1 FILLER_0_11_160 ();
 FILLCELL_X2 FILLER_0_11_167 ();
 FILLCELL_X16 FILLER_0_11_183 ();
 FILLCELL_X4 FILLER_0_11_199 ();
 FILLCELL_X2 FILLER_0_11_213 ();
 FILLCELL_X1 FILLER_0_11_215 ();
 FILLCELL_X1 FILLER_0_11_228 ();
 FILLCELL_X8 FILLER_0_11_243 ();
 FILLCELL_X4 FILLER_0_11_251 ();
 FILLCELL_X4 FILLER_0_11_263 ();
 FILLCELL_X1 FILLER_0_11_267 ();
 FILLCELL_X2 FILLER_0_11_270 ();
 FILLCELL_X4 FILLER_0_11_276 ();
 FILLCELL_X1 FILLER_0_11_280 ();
 FILLCELL_X4 FILLER_0_11_283 ();
 FILLCELL_X2 FILLER_0_11_287 ();
 FILLCELL_X1 FILLER_0_11_289 ();
 FILLCELL_X1 FILLER_0_11_345 ();
 FILLCELL_X1 FILLER_0_11_370 ();
 FILLCELL_X8 FILLER_0_11_380 ();
 FILLCELL_X2 FILLER_0_12_1 ();
 FILLCELL_X2 FILLER_0_12_7 ();
 FILLCELL_X1 FILLER_0_12_9 ();
 FILLCELL_X1 FILLER_0_12_13 ();
 FILLCELL_X2 FILLER_0_12_18 ();
 FILLCELL_X1 FILLER_0_12_20 ();
 FILLCELL_X1 FILLER_0_12_25 ();
 FILLCELL_X2 FILLER_0_12_48 ();
 FILLCELL_X1 FILLER_0_12_58 ();
 FILLCELL_X8 FILLER_0_12_63 ();
 FILLCELL_X4 FILLER_0_12_84 ();
 FILLCELL_X1 FILLER_0_12_88 ();
 FILLCELL_X1 FILLER_0_12_112 ();
 FILLCELL_X1 FILLER_0_12_116 ();
 FILLCELL_X2 FILLER_0_12_123 ();
 FILLCELL_X1 FILLER_0_12_125 ();
 FILLCELL_X4 FILLER_0_12_132 ();
 FILLCELL_X4 FILLER_0_12_139 ();
 FILLCELL_X1 FILLER_0_12_143 ();
 FILLCELL_X8 FILLER_0_12_160 ();
 FILLCELL_X2 FILLER_0_12_168 ();
 FILLCELL_X1 FILLER_0_12_170 ();
 FILLCELL_X1 FILLER_0_12_217 ();
 FILLCELL_X2 FILLER_0_12_224 ();
 FILLCELL_X2 FILLER_0_12_230 ();
 FILLCELL_X2 FILLER_0_12_238 ();
 FILLCELL_X4 FILLER_0_12_244 ();
 FILLCELL_X2 FILLER_0_12_248 ();
 FILLCELL_X1 FILLER_0_12_250 ();
 FILLCELL_X1 FILLER_0_12_266 ();
 FILLCELL_X2 FILLER_0_12_284 ();
 FILLCELL_X1 FILLER_0_12_289 ();
 FILLCELL_X2 FILLER_0_12_296 ();
 FILLCELL_X1 FILLER_0_12_307 ();
 FILLCELL_X1 FILLER_0_12_321 ();
 FILLCELL_X2 FILLER_0_12_325 ();
 FILLCELL_X2 FILLER_0_12_330 ();
 FILLCELL_X2 FILLER_0_12_338 ();
 FILLCELL_X1 FILLER_0_12_349 ();
 FILLCELL_X2 FILLER_0_12_378 ();
 FILLCELL_X4 FILLER_0_12_384 ();
 FILLCELL_X2 FILLER_0_13_1 ();
 FILLCELL_X1 FILLER_0_13_10 ();
 FILLCELL_X1 FILLER_0_13_17 ();
 FILLCELL_X1 FILLER_0_13_21 ();
 FILLCELL_X2 FILLER_0_13_27 ();
 FILLCELL_X4 FILLER_0_13_38 ();
 FILLCELL_X2 FILLER_0_13_42 ();
 FILLCELL_X1 FILLER_0_13_44 ();
 FILLCELL_X4 FILLER_0_13_58 ();
 FILLCELL_X2 FILLER_0_13_62 ();
 FILLCELL_X1 FILLER_0_13_64 ();
 FILLCELL_X1 FILLER_0_13_74 ();
 FILLCELL_X1 FILLER_0_13_78 ();
 FILLCELL_X1 FILLER_0_13_85 ();
 FILLCELL_X1 FILLER_0_13_92 ();
 FILLCELL_X1 FILLER_0_13_96 ();
 FILLCELL_X1 FILLER_0_13_101 ();
 FILLCELL_X1 FILLER_0_13_106 ();
 FILLCELL_X2 FILLER_0_13_113 ();
 FILLCELL_X1 FILLER_0_13_119 ();
 FILLCELL_X2 FILLER_0_13_122 ();
 FILLCELL_X1 FILLER_0_13_124 ();
 FILLCELL_X2 FILLER_0_13_131 ();
 FILLCELL_X1 FILLER_0_13_144 ();
 FILLCELL_X1 FILLER_0_13_151 ();
 FILLCELL_X1 FILLER_0_13_155 ();
 FILLCELL_X1 FILLER_0_13_160 ();
 FILLCELL_X1 FILLER_0_13_167 ();
 FILLCELL_X4 FILLER_0_13_171 ();
 FILLCELL_X2 FILLER_0_13_175 ();
 FILLCELL_X1 FILLER_0_13_177 ();
 FILLCELL_X4 FILLER_0_13_185 ();
 FILLCELL_X8 FILLER_0_13_211 ();
 FILLCELL_X4 FILLER_0_13_219 ();
 FILLCELL_X1 FILLER_0_13_223 ();
 FILLCELL_X4 FILLER_0_13_230 ();
 FILLCELL_X8 FILLER_0_13_237 ();
 FILLCELL_X4 FILLER_0_13_245 ();
 FILLCELL_X2 FILLER_0_13_249 ();
 FILLCELL_X2 FILLER_0_13_288 ();
 FILLCELL_X1 FILLER_0_13_290 ();
 FILLCELL_X2 FILLER_0_13_307 ();
 FILLCELL_X2 FILLER_0_13_320 ();
 FILLCELL_X1 FILLER_0_13_322 ();
 FILLCELL_X2 FILLER_0_13_340 ();
 FILLCELL_X4 FILLER_0_13_346 ();
 FILLCELL_X1 FILLER_0_13_357 ();
 FILLCELL_X1 FILLER_0_13_361 ();
 FILLCELL_X1 FILLER_0_13_383 ();
 FILLCELL_X4 FILLER_0_14_13 ();
 FILLCELL_X1 FILLER_0_14_17 ();
 FILLCELL_X2 FILLER_0_14_38 ();
 FILLCELL_X1 FILLER_0_14_40 ();
 FILLCELL_X2 FILLER_0_14_47 ();
 FILLCELL_X1 FILLER_0_14_52 ();
 FILLCELL_X1 FILLER_0_14_62 ();
 FILLCELL_X1 FILLER_0_14_76 ();
 FILLCELL_X2 FILLER_0_14_83 ();
 FILLCELL_X1 FILLER_0_14_85 ();
 FILLCELL_X1 FILLER_0_14_90 ();
 FILLCELL_X1 FILLER_0_14_109 ();
 FILLCELL_X1 FILLER_0_14_114 ();
 FILLCELL_X1 FILLER_0_14_130 ();
 FILLCELL_X1 FILLER_0_14_137 ();
 FILLCELL_X1 FILLER_0_14_163 ();
 FILLCELL_X1 FILLER_0_14_170 ();
 FILLCELL_X1 FILLER_0_14_173 ();
 FILLCELL_X1 FILLER_0_14_180 ();
 FILLCELL_X4 FILLER_0_14_185 ();
 FILLCELL_X1 FILLER_0_14_189 ();
 FILLCELL_X8 FILLER_0_14_199 ();
 FILLCELL_X4 FILLER_0_14_242 ();
 FILLCELL_X2 FILLER_0_14_246 ();
 FILLCELL_X2 FILLER_0_14_265 ();
 FILLCELL_X4 FILLER_0_14_305 ();
 FILLCELL_X1 FILLER_0_14_330 ();
 FILLCELL_X1 FILLER_0_14_337 ();
 FILLCELL_X1 FILLER_0_14_344 ();
 FILLCELL_X2 FILLER_0_14_349 ();
 FILLCELL_X2 FILLER_0_14_354 ();
 FILLCELL_X1 FILLER_0_14_356 ();
 FILLCELL_X1 FILLER_0_14_361 ();
 FILLCELL_X1 FILLER_0_14_365 ();
 FILLCELL_X4 FILLER_0_14_383 ();
 FILLCELL_X1 FILLER_0_14_387 ();
 FILLCELL_X8 FILLER_0_15_11 ();
 FILLCELL_X1 FILLER_0_15_29 ();
 FILLCELL_X4 FILLER_0_15_39 ();
 FILLCELL_X1 FILLER_0_15_43 ();
 FILLCELL_X2 FILLER_0_15_50 ();
 FILLCELL_X4 FILLER_0_15_59 ();
 FILLCELL_X2 FILLER_0_15_69 ();
 FILLCELL_X1 FILLER_0_15_71 ();
 FILLCELL_X2 FILLER_0_15_76 ();
 FILLCELL_X1 FILLER_0_15_78 ();
 FILLCELL_X1 FILLER_0_15_107 ();
 FILLCELL_X4 FILLER_0_15_114 ();
 FILLCELL_X2 FILLER_0_15_118 ();
 FILLCELL_X2 FILLER_0_15_134 ();
 FILLCELL_X1 FILLER_0_15_136 ();
 FILLCELL_X1 FILLER_0_15_181 ();
 FILLCELL_X1 FILLER_0_15_204 ();
 FILLCELL_X2 FILLER_0_15_220 ();
 FILLCELL_X2 FILLER_0_15_226 ();
 FILLCELL_X1 FILLER_0_15_251 ();
 FILLCELL_X2 FILLER_0_15_267 ();
 FILLCELL_X1 FILLER_0_15_269 ();
 FILLCELL_X4 FILLER_0_15_278 ();
 FILLCELL_X1 FILLER_0_15_282 ();
 FILLCELL_X1 FILLER_0_15_326 ();
 FILLCELL_X2 FILLER_0_15_351 ();
 FILLCELL_X1 FILLER_0_15_381 ();
 FILLCELL_X2 FILLER_0_15_386 ();
 FILLCELL_X8 FILLER_0_16_9 ();
 FILLCELL_X4 FILLER_0_16_17 ();
 FILLCELL_X2 FILLER_0_16_21 ();
 FILLCELL_X1 FILLER_0_16_23 ();
 FILLCELL_X1 FILLER_0_16_52 ();
 FILLCELL_X1 FILLER_0_16_59 ();
 FILLCELL_X1 FILLER_0_16_70 ();
 FILLCELL_X2 FILLER_0_16_87 ();
 FILLCELL_X2 FILLER_0_16_90 ();
 FILLCELL_X2 FILLER_0_16_111 ();
 FILLCELL_X1 FILLER_0_16_113 ();
 FILLCELL_X1 FILLER_0_16_118 ();
 FILLCELL_X2 FILLER_0_16_159 ();
 FILLCELL_X1 FILLER_0_16_167 ();
 FILLCELL_X2 FILLER_0_16_178 ();
 FILLCELL_X1 FILLER_0_16_211 ();
 FILLCELL_X1 FILLER_0_16_215 ();
 FILLCELL_X1 FILLER_0_16_225 ();
 FILLCELL_X1 FILLER_0_16_238 ();
 FILLCELL_X2 FILLER_0_16_242 ();
 FILLCELL_X1 FILLER_0_16_244 ();
 FILLCELL_X8 FILLER_0_16_255 ();
 FILLCELL_X4 FILLER_0_16_263 ();
 FILLCELL_X4 FILLER_0_16_268 ();
 FILLCELL_X2 FILLER_0_16_272 ();
 FILLCELL_X1 FILLER_0_16_274 ();
 FILLCELL_X1 FILLER_0_16_281 ();
 FILLCELL_X4 FILLER_0_16_288 ();
 FILLCELL_X2 FILLER_0_16_295 ();
 FILLCELL_X4 FILLER_0_16_300 ();
 FILLCELL_X2 FILLER_0_16_304 ();
 FILLCELL_X4 FILLER_0_16_316 ();
 FILLCELL_X2 FILLER_0_16_341 ();
 FILLCELL_X1 FILLER_0_16_363 ();
 FILLCELL_X4 FILLER_0_16_383 ();
 FILLCELL_X1 FILLER_0_16_387 ();
 FILLCELL_X2 FILLER_0_17_1 ();
 FILLCELL_X8 FILLER_0_17_23 ();
 FILLCELL_X1 FILLER_0_17_37 ();
 FILLCELL_X1 FILLER_0_17_44 ();
 FILLCELL_X2 FILLER_0_17_61 ();
 FILLCELL_X2 FILLER_0_17_76 ();
 FILLCELL_X1 FILLER_0_17_87 ();
 FILLCELL_X1 FILLER_0_17_91 ();
 FILLCELL_X1 FILLER_0_17_99 ();
 FILLCELL_X4 FILLER_0_17_112 ();
 FILLCELL_X1 FILLER_0_17_120 ();
 FILLCELL_X1 FILLER_0_17_130 ();
 FILLCELL_X2 FILLER_0_17_137 ();
 FILLCELL_X1 FILLER_0_17_151 ();
 FILLCELL_X1 FILLER_0_17_156 ();
 FILLCELL_X1 FILLER_0_17_169 ();
 FILLCELL_X1 FILLER_0_17_179 ();
 FILLCELL_X2 FILLER_0_17_193 ();
 FILLCELL_X1 FILLER_0_17_195 ();
 FILLCELL_X4 FILLER_0_17_207 ();
 FILLCELL_X1 FILLER_0_17_237 ();
 FILLCELL_X1 FILLER_0_17_245 ();
 FILLCELL_X4 FILLER_0_17_253 ();
 FILLCELL_X8 FILLER_0_17_274 ();
 FILLCELL_X4 FILLER_0_17_282 ();
 FILLCELL_X1 FILLER_0_17_312 ();
 FILLCELL_X1 FILLER_0_17_320 ();
 FILLCELL_X1 FILLER_0_17_324 ();
 FILLCELL_X1 FILLER_0_17_329 ();
 FILLCELL_X2 FILLER_0_17_333 ();
 FILLCELL_X1 FILLER_0_17_335 ();
 FILLCELL_X4 FILLER_0_17_350 ();
 FILLCELL_X2 FILLER_0_17_354 ();
 FILLCELL_X4 FILLER_0_17_363 ();
 FILLCELL_X1 FILLER_0_17_367 ();
 FILLCELL_X1 FILLER_0_18_22 ();
 FILLCELL_X1 FILLER_0_18_32 ();
 FILLCELL_X1 FILLER_0_18_47 ();
 FILLCELL_X1 FILLER_0_18_54 ();
 FILLCELL_X2 FILLER_0_18_68 ();
 FILLCELL_X2 FILLER_0_18_76 ();
 FILLCELL_X1 FILLER_0_18_78 ();
 FILLCELL_X2 FILLER_0_18_85 ();
 FILLCELL_X2 FILLER_0_18_136 ();
 FILLCELL_X2 FILLER_0_18_153 ();
 FILLCELL_X1 FILLER_0_18_155 ();
 FILLCELL_X2 FILLER_0_18_165 ();
 FILLCELL_X1 FILLER_0_18_174 ();
 FILLCELL_X4 FILLER_0_18_177 ();
 FILLCELL_X2 FILLER_0_18_181 ();
 FILLCELL_X1 FILLER_0_18_185 ();
 FILLCELL_X1 FILLER_0_18_192 ();
 FILLCELL_X2 FILLER_0_18_199 ();
 FILLCELL_X1 FILLER_0_18_204 ();
 FILLCELL_X2 FILLER_0_18_209 ();
 FILLCELL_X4 FILLER_0_18_220 ();
 FILLCELL_X1 FILLER_0_18_224 ();
 FILLCELL_X4 FILLER_0_18_234 ();
 FILLCELL_X2 FILLER_0_18_238 ();
 FILLCELL_X4 FILLER_0_18_268 ();
 FILLCELL_X1 FILLER_0_18_285 ();
 FILLCELL_X1 FILLER_0_18_310 ();
 FILLCELL_X2 FILLER_0_18_317 ();
 FILLCELL_X8 FILLER_0_18_325 ();
 FILLCELL_X4 FILLER_0_18_333 ();
 FILLCELL_X2 FILLER_0_18_337 ();
 FILLCELL_X1 FILLER_0_18_339 ();
 FILLCELL_X2 FILLER_0_18_367 ();
 FILLCELL_X2 FILLER_0_18_386 ();
 FILLCELL_X4 FILLER_0_19_1 ();
 FILLCELL_X2 FILLER_0_19_5 ();
 FILLCELL_X4 FILLER_0_19_19 ();
 FILLCELL_X2 FILLER_0_19_23 ();
 FILLCELL_X1 FILLER_0_19_25 ();
 FILLCELL_X1 FILLER_0_19_32 ();
 FILLCELL_X1 FILLER_0_19_54 ();
 FILLCELL_X2 FILLER_0_19_84 ();
 FILLCELL_X1 FILLER_0_19_86 ();
 FILLCELL_X4 FILLER_0_19_93 ();
 FILLCELL_X2 FILLER_0_19_97 ();
 FILLCELL_X1 FILLER_0_19_99 ();
 FILLCELL_X2 FILLER_0_19_143 ();
 FILLCELL_X1 FILLER_0_19_156 ();
 FILLCELL_X2 FILLER_0_19_176 ();
 FILLCELL_X1 FILLER_0_19_206 ();
 FILLCELL_X1 FILLER_0_19_212 ();
 FILLCELL_X4 FILLER_0_19_221 ();
 FILLCELL_X2 FILLER_0_19_225 ();
 FILLCELL_X2 FILLER_0_19_244 ();
 FILLCELL_X2 FILLER_0_19_249 ();
 FILLCELL_X2 FILLER_0_19_257 ();
 FILLCELL_X8 FILLER_0_19_269 ();
 FILLCELL_X2 FILLER_0_19_277 ();
 FILLCELL_X2 FILLER_0_19_292 ();
 FILLCELL_X1 FILLER_0_19_294 ();
 FILLCELL_X1 FILLER_0_19_316 ();
 FILLCELL_X2 FILLER_0_19_330 ();
 FILLCELL_X1 FILLER_0_19_332 ();
 FILLCELL_X2 FILLER_0_19_336 ();
 FILLCELL_X4 FILLER_0_19_357 ();
 FILLCELL_X2 FILLER_0_19_361 ();
 FILLCELL_X2 FILLER_0_19_382 ();
 FILLCELL_X1 FILLER_0_19_387 ();
 FILLCELL_X2 FILLER_0_20_1 ();
 FILLCELL_X2 FILLER_0_20_31 ();
 FILLCELL_X2 FILLER_0_20_37 ();
 FILLCELL_X1 FILLER_0_20_59 ();
 FILLCELL_X1 FILLER_0_20_63 ();
 FILLCELL_X1 FILLER_0_20_68 ();
 FILLCELL_X1 FILLER_0_20_75 ();
 FILLCELL_X1 FILLER_0_20_79 ();
 FILLCELL_X2 FILLER_0_20_84 ();
 FILLCELL_X1 FILLER_0_20_90 ();
 FILLCELL_X2 FILLER_0_20_97 ();
 FILLCELL_X1 FILLER_0_20_99 ();
 FILLCELL_X1 FILLER_0_20_163 ();
 FILLCELL_X4 FILLER_0_20_174 ();
 FILLCELL_X1 FILLER_0_20_184 ();
 FILLCELL_X2 FILLER_0_20_187 ();
 FILLCELL_X1 FILLER_0_20_195 ();
 FILLCELL_X2 FILLER_0_20_202 ();
 FILLCELL_X4 FILLER_0_20_233 ();
 FILLCELL_X2 FILLER_0_20_237 ();
 FILLCELL_X1 FILLER_0_20_245 ();
 FILLCELL_X1 FILLER_0_20_249 ();
 FILLCELL_X1 FILLER_0_20_257 ();
 FILLCELL_X1 FILLER_0_20_260 ();
 FILLCELL_X2 FILLER_0_20_268 ();
 FILLCELL_X2 FILLER_0_20_273 ();
 FILLCELL_X1 FILLER_0_20_275 ();
 FILLCELL_X8 FILLER_0_20_278 ();
 FILLCELL_X2 FILLER_0_20_292 ();
 FILLCELL_X1 FILLER_0_20_300 ();
 FILLCELL_X1 FILLER_0_20_307 ();
 FILLCELL_X4 FILLER_0_20_359 ();
 FILLCELL_X2 FILLER_0_20_363 ();
 FILLCELL_X2 FILLER_0_20_382 ();
 FILLCELL_X2 FILLER_0_21_1 ();
 FILLCELL_X4 FILLER_0_21_10 ();
 FILLCELL_X2 FILLER_0_21_14 ();
 FILLCELL_X1 FILLER_0_21_16 ();
 FILLCELL_X2 FILLER_0_21_25 ();
 FILLCELL_X1 FILLER_0_21_27 ();
 FILLCELL_X1 FILLER_0_21_31 ();
 FILLCELL_X2 FILLER_0_21_62 ();
 FILLCELL_X2 FILLER_0_21_67 ();
 FILLCELL_X1 FILLER_0_21_69 ();
 FILLCELL_X2 FILLER_0_21_92 ();
 FILLCELL_X1 FILLER_0_21_98 ();
 FILLCELL_X1 FILLER_0_21_102 ();
 FILLCELL_X1 FILLER_0_21_122 ();
 FILLCELL_X4 FILLER_0_21_129 ();
 FILLCELL_X1 FILLER_0_21_150 ();
 FILLCELL_X1 FILLER_0_21_171 ();
 FILLCELL_X1 FILLER_0_21_191 ();
 FILLCELL_X8 FILLER_0_21_196 ();
 FILLCELL_X2 FILLER_0_21_204 ();
 FILLCELL_X1 FILLER_0_21_206 ();
 FILLCELL_X2 FILLER_0_21_216 ();
 FILLCELL_X1 FILLER_0_21_232 ();
 FILLCELL_X2 FILLER_0_21_262 ();
 FILLCELL_X1 FILLER_0_21_264 ();
 FILLCELL_X2 FILLER_0_21_285 ();
 FILLCELL_X1 FILLER_0_21_287 ();
 FILLCELL_X8 FILLER_0_21_304 ();
 FILLCELL_X8 FILLER_0_21_331 ();
 FILLCELL_X2 FILLER_0_21_339 ();
 FILLCELL_X1 FILLER_0_21_341 ();
 FILLCELL_X1 FILLER_0_21_379 ();
 FILLCELL_X2 FILLER_0_21_386 ();
 FILLCELL_X1 FILLER_0_22_13 ();
 FILLCELL_X2 FILLER_0_22_17 ();
 FILLCELL_X2 FILLER_0_22_25 ();
 FILLCELL_X2 FILLER_0_22_33 ();
 FILLCELL_X4 FILLER_0_22_41 ();
 FILLCELL_X1 FILLER_0_22_69 ();
 FILLCELL_X4 FILLER_0_22_73 ();
 FILLCELL_X2 FILLER_0_22_80 ();
 FILLCELL_X1 FILLER_0_22_90 ();
 FILLCELL_X1 FILLER_0_22_97 ();
 FILLCELL_X1 FILLER_0_22_102 ();
 FILLCELL_X2 FILLER_0_22_121 ();
 FILLCELL_X1 FILLER_0_22_129 ();
 FILLCELL_X1 FILLER_0_22_136 ();
 FILLCELL_X2 FILLER_0_22_142 ();
 FILLCELL_X1 FILLER_0_22_150 ();
 FILLCELL_X1 FILLER_0_22_154 ();
 FILLCELL_X1 FILLER_0_22_158 ();
 FILLCELL_X1 FILLER_0_22_161 ();
 FILLCELL_X1 FILLER_0_22_168 ();
 FILLCELL_X2 FILLER_0_22_171 ();
 FILLCELL_X8 FILLER_0_22_189 ();
 FILLCELL_X4 FILLER_0_22_197 ();
 FILLCELL_X2 FILLER_0_22_231 ();
 FILLCELL_X1 FILLER_0_22_233 ();
 FILLCELL_X4 FILLER_0_22_247 ();
 FILLCELL_X2 FILLER_0_22_251 ();
 FILLCELL_X4 FILLER_0_22_262 ();
 FILLCELL_X1 FILLER_0_22_266 ();
 FILLCELL_X4 FILLER_0_22_268 ();
 FILLCELL_X1 FILLER_0_22_287 ();
 FILLCELL_X4 FILLER_0_22_311 ();
 FILLCELL_X4 FILLER_0_22_328 ();
 FILLCELL_X2 FILLER_0_22_332 ();
 FILLCELL_X1 FILLER_0_22_344 ();
 FILLCELL_X2 FILLER_0_22_380 ();
 FILLCELL_X1 FILLER_0_23_1 ();
 FILLCELL_X1 FILLER_0_23_8 ();
 FILLCELL_X1 FILLER_0_23_12 ();
 FILLCELL_X2 FILLER_0_23_19 ();
 FILLCELL_X2 FILLER_0_23_27 ();
 FILLCELL_X2 FILLER_0_23_35 ();
 FILLCELL_X1 FILLER_0_23_37 ();
 FILLCELL_X1 FILLER_0_23_43 ();
 FILLCELL_X8 FILLER_0_23_50 ();
 FILLCELL_X2 FILLER_0_23_58 ();
 FILLCELL_X4 FILLER_0_23_66 ();
 FILLCELL_X1 FILLER_0_23_70 ();
 FILLCELL_X1 FILLER_0_23_75 ();
 FILLCELL_X1 FILLER_0_23_89 ();
 FILLCELL_X1 FILLER_0_23_96 ();
 FILLCELL_X1 FILLER_0_23_103 ();
 FILLCELL_X1 FILLER_0_23_120 ();
 FILLCELL_X1 FILLER_0_23_127 ();
 FILLCELL_X1 FILLER_0_23_133 ();
 FILLCELL_X2 FILLER_0_23_140 ();
 FILLCELL_X1 FILLER_0_23_142 ();
 FILLCELL_X4 FILLER_0_23_149 ();
 FILLCELL_X2 FILLER_0_23_153 ();
 FILLCELL_X1 FILLER_0_23_155 ();
 FILLCELL_X2 FILLER_0_23_169 ();
 FILLCELL_X1 FILLER_0_23_171 ();
 FILLCELL_X2 FILLER_0_23_179 ();
 FILLCELL_X8 FILLER_0_23_185 ();
 FILLCELL_X4 FILLER_0_23_193 ();
 FILLCELL_X2 FILLER_0_23_197 ();
 FILLCELL_X4 FILLER_0_23_207 ();
 FILLCELL_X4 FILLER_0_23_216 ();
 FILLCELL_X4 FILLER_0_23_231 ();
 FILLCELL_X1 FILLER_0_23_235 ();
 FILLCELL_X2 FILLER_0_23_250 ();
 FILLCELL_X2 FILLER_0_23_255 ();
 FILLCELL_X1 FILLER_0_23_261 ();
 FILLCELL_X2 FILLER_0_23_268 ();
 FILLCELL_X1 FILLER_0_23_270 ();
 FILLCELL_X2 FILLER_0_23_277 ();
 FILLCELL_X2 FILLER_0_23_289 ();
 FILLCELL_X4 FILLER_0_23_297 ();
 FILLCELL_X2 FILLER_0_23_301 ();
 FILLCELL_X1 FILLER_0_23_303 ();
 FILLCELL_X1 FILLER_0_23_314 ();
 FILLCELL_X4 FILLER_0_23_324 ();
 FILLCELL_X2 FILLER_0_23_328 ();
 FILLCELL_X1 FILLER_0_23_330 ();
 FILLCELL_X1 FILLER_0_23_349 ();
 FILLCELL_X1 FILLER_0_23_379 ();
 FILLCELL_X4 FILLER_0_23_384 ();
 FILLCELL_X8 FILLER_0_24_1 ();
 FILLCELL_X1 FILLER_0_24_9 ();
 FILLCELL_X2 FILLER_0_24_22 ();
 FILLCELL_X1 FILLER_0_24_30 ();
 FILLCELL_X2 FILLER_0_24_44 ();
 FILLCELL_X1 FILLER_0_24_50 ();
 FILLCELL_X2 FILLER_0_24_86 ();
 FILLCELL_X1 FILLER_0_24_88 ();
 FILLCELL_X2 FILLER_0_24_90 ();
 FILLCELL_X1 FILLER_0_24_92 ();
 FILLCELL_X2 FILLER_0_24_96 ();
 FILLCELL_X1 FILLER_0_24_98 ();
 FILLCELL_X2 FILLER_0_24_112 ();
 FILLCELL_X1 FILLER_0_24_114 ();
 FILLCELL_X4 FILLER_0_24_130 ();
 FILLCELL_X1 FILLER_0_24_134 ();
 FILLCELL_X2 FILLER_0_24_139 ();
 FILLCELL_X8 FILLER_0_24_150 ();
 FILLCELL_X2 FILLER_0_24_158 ();
 FILLCELL_X8 FILLER_0_24_170 ();
 FILLCELL_X1 FILLER_0_24_187 ();
 FILLCELL_X1 FILLER_0_24_194 ();
 FILLCELL_X1 FILLER_0_24_199 ();
 FILLCELL_X1 FILLER_0_24_204 ();
 FILLCELL_X2 FILLER_0_24_208 ();
 FILLCELL_X8 FILLER_0_24_213 ();
 FILLCELL_X4 FILLER_0_24_221 ();
 FILLCELL_X1 FILLER_0_24_225 ();
 FILLCELL_X2 FILLER_0_24_241 ();
 FILLCELL_X1 FILLER_0_24_249 ();
 FILLCELL_X8 FILLER_0_24_268 ();
 FILLCELL_X2 FILLER_0_24_276 ();
 FILLCELL_X1 FILLER_0_24_297 ();
 FILLCELL_X1 FILLER_0_24_301 ();
 FILLCELL_X1 FILLER_0_24_308 ();
 FILLCELL_X1 FILLER_0_24_312 ();
 FILLCELL_X1 FILLER_0_24_317 ();
 FILLCELL_X1 FILLER_0_24_321 ();
 FILLCELL_X1 FILLER_0_24_326 ();
 FILLCELL_X1 FILLER_0_24_332 ();
 FILLCELL_X1 FILLER_0_24_354 ();
 FILLCELL_X1 FILLER_0_24_358 ();
 FILLCELL_X2 FILLER_0_24_361 ();
 FILLCELL_X2 FILLER_0_24_369 ();
 FILLCELL_X4 FILLER_0_25_1 ();
 FILLCELL_X2 FILLER_0_25_5 ();
 FILLCELL_X1 FILLER_0_25_7 ();
 FILLCELL_X2 FILLER_0_25_24 ();
 FILLCELL_X2 FILLER_0_25_48 ();
 FILLCELL_X4 FILLER_0_25_53 ();
 FILLCELL_X1 FILLER_0_25_57 ();
 FILLCELL_X1 FILLER_0_25_65 ();
 FILLCELL_X1 FILLER_0_25_72 ();
 FILLCELL_X8 FILLER_0_25_86 ();
 FILLCELL_X4 FILLER_0_25_94 ();
 FILLCELL_X2 FILLER_0_25_98 ();
 FILLCELL_X2 FILLER_0_25_121 ();
 FILLCELL_X2 FILLER_0_25_127 ();
 FILLCELL_X1 FILLER_0_25_129 ();
 FILLCELL_X2 FILLER_0_25_136 ();
 FILLCELL_X2 FILLER_0_25_147 ();
 FILLCELL_X1 FILLER_0_25_153 ();
 FILLCELL_X4 FILLER_0_25_166 ();
 FILLCELL_X2 FILLER_0_25_172 ();
 FILLCELL_X1 FILLER_0_25_174 ();
 FILLCELL_X1 FILLER_0_25_179 ();
 FILLCELL_X1 FILLER_0_25_186 ();
 FILLCELL_X1 FILLER_0_25_197 ();
 FILLCELL_X4 FILLER_0_25_202 ();
 FILLCELL_X1 FILLER_0_25_206 ();
 FILLCELL_X4 FILLER_0_25_224 ();
 FILLCELL_X1 FILLER_0_25_228 ();
 FILLCELL_X2 FILLER_0_25_245 ();
 FILLCELL_X1 FILLER_0_25_247 ();
 FILLCELL_X4 FILLER_0_25_254 ();
 FILLCELL_X2 FILLER_0_25_258 ();
 FILLCELL_X1 FILLER_0_25_260 ();
 FILLCELL_X1 FILLER_0_25_290 ();
 FILLCELL_X1 FILLER_0_25_298 ();
 FILLCELL_X1 FILLER_0_25_307 ();
 FILLCELL_X4 FILLER_0_25_314 ();
 FILLCELL_X1 FILLER_0_25_318 ();
 FILLCELL_X2 FILLER_0_25_347 ();
 FILLCELL_X8 FILLER_0_25_377 ();
 FILLCELL_X2 FILLER_0_25_385 ();
 FILLCELL_X1 FILLER_0_25_387 ();
 FILLCELL_X2 FILLER_0_26_38 ();
 FILLCELL_X1 FILLER_0_26_55 ();
 FILLCELL_X1 FILLER_0_26_62 ();
 FILLCELL_X1 FILLER_0_26_72 ();
 FILLCELL_X4 FILLER_0_26_75 ();
 FILLCELL_X4 FILLER_0_26_85 ();
 FILLCELL_X1 FILLER_0_26_90 ();
 FILLCELL_X1 FILLER_0_26_100 ();
 FILLCELL_X1 FILLER_0_26_105 ();
 FILLCELL_X1 FILLER_0_26_115 ();
 FILLCELL_X1 FILLER_0_26_122 ();
 FILLCELL_X1 FILLER_0_26_127 ();
 FILLCELL_X8 FILLER_0_26_133 ();
 FILLCELL_X4 FILLER_0_26_141 ();
 FILLCELL_X2 FILLER_0_26_145 ();
 FILLCELL_X2 FILLER_0_26_169 ();
 FILLCELL_X1 FILLER_0_26_171 ();
 FILLCELL_X2 FILLER_0_26_179 ();
 FILLCELL_X1 FILLER_0_26_185 ();
 FILLCELL_X2 FILLER_0_26_193 ();
 FILLCELL_X1 FILLER_0_26_195 ();
 FILLCELL_X1 FILLER_0_26_203 ();
 FILLCELL_X8 FILLER_0_26_210 ();
 FILLCELL_X1 FILLER_0_26_218 ();
 FILLCELL_X2 FILLER_0_26_231 ();
 FILLCELL_X1 FILLER_0_26_233 ();
 FILLCELL_X2 FILLER_0_26_240 ();
 FILLCELL_X2 FILLER_0_26_265 ();
 FILLCELL_X4 FILLER_0_26_268 ();
 FILLCELL_X2 FILLER_0_26_272 ();
 FILLCELL_X1 FILLER_0_26_274 ();
 FILLCELL_X2 FILLER_0_26_290 ();
 FILLCELL_X2 FILLER_0_26_301 ();
 FILLCELL_X2 FILLER_0_26_338 ();
 FILLCELL_X2 FILLER_0_26_358 ();
 FILLCELL_X2 FILLER_0_26_366 ();
 FILLCELL_X1 FILLER_0_27_10 ();
 FILLCELL_X2 FILLER_0_27_30 ();
 FILLCELL_X8 FILLER_0_27_78 ();
 FILLCELL_X2 FILLER_0_27_86 ();
 FILLCELL_X1 FILLER_0_27_103 ();
 FILLCELL_X1 FILLER_0_27_120 ();
 FILLCELL_X8 FILLER_0_27_134 ();
 FILLCELL_X4 FILLER_0_27_142 ();
 FILLCELL_X1 FILLER_0_27_146 ();
 FILLCELL_X2 FILLER_0_27_160 ();
 FILLCELL_X1 FILLER_0_27_162 ();
 FILLCELL_X1 FILLER_0_27_171 ();
 FILLCELL_X4 FILLER_0_27_179 ();
 FILLCELL_X2 FILLER_0_27_193 ();
 FILLCELL_X1 FILLER_0_27_195 ();
 FILLCELL_X1 FILLER_0_27_202 ();
 FILLCELL_X8 FILLER_0_27_207 ();
 FILLCELL_X4 FILLER_0_27_215 ();
 FILLCELL_X2 FILLER_0_27_219 ();
 FILLCELL_X1 FILLER_0_27_227 ();
 FILLCELL_X1 FILLER_0_27_232 ();
 FILLCELL_X1 FILLER_0_27_241 ();
 FILLCELL_X4 FILLER_0_27_245 ();
 FILLCELL_X4 FILLER_0_27_259 ();
 FILLCELL_X1 FILLER_0_27_282 ();
 FILLCELL_X2 FILLER_0_27_296 ();
 FILLCELL_X4 FILLER_0_27_308 ();
 FILLCELL_X1 FILLER_0_27_312 ();
 FILLCELL_X2 FILLER_0_27_316 ();
 FILLCELL_X1 FILLER_0_27_324 ();
 FILLCELL_X8 FILLER_0_27_334 ();
 FILLCELL_X2 FILLER_0_27_342 ();
 FILLCELL_X1 FILLER_0_27_344 ();
 FILLCELL_X1 FILLER_0_27_352 ();
 FILLCELL_X1 FILLER_0_27_374 ();
 FILLCELL_X4 FILLER_0_27_381 ();
 FILLCELL_X2 FILLER_0_27_385 ();
 FILLCELL_X1 FILLER_0_27_387 ();
 FILLCELL_X4 FILLER_0_28_1 ();
 FILLCELL_X1 FILLER_0_28_5 ();
 FILLCELL_X2 FILLER_0_28_12 ();
 FILLCELL_X1 FILLER_0_28_20 ();
 FILLCELL_X2 FILLER_0_28_24 ();
 FILLCELL_X1 FILLER_0_28_29 ();
 FILLCELL_X2 FILLER_0_28_43 ();
 FILLCELL_X1 FILLER_0_28_45 ();
 FILLCELL_X2 FILLER_0_28_52 ();
 FILLCELL_X1 FILLER_0_28_82 ();
 FILLCELL_X4 FILLER_0_28_94 ();
 FILLCELL_X1 FILLER_0_28_98 ();
 FILLCELL_X2 FILLER_0_28_133 ();
 FILLCELL_X8 FILLER_0_28_141 ();
 FILLCELL_X1 FILLER_0_28_149 ();
 FILLCELL_X1 FILLER_0_28_167 ();
 FILLCELL_X2 FILLER_0_28_174 ();
 FILLCELL_X2 FILLER_0_28_179 ();
 FILLCELL_X1 FILLER_0_28_190 ();
 FILLCELL_X1 FILLER_0_28_223 ();
 FILLCELL_X1 FILLER_0_28_250 ();
 FILLCELL_X4 FILLER_0_28_254 ();
 FILLCELL_X2 FILLER_0_28_258 ();
 FILLCELL_X1 FILLER_0_28_266 ();
 FILLCELL_X1 FILLER_0_28_272 ();
 FILLCELL_X1 FILLER_0_28_277 ();
 FILLCELL_X2 FILLER_0_28_282 ();
 FILLCELL_X2 FILLER_0_28_290 ();
 FILLCELL_X4 FILLER_0_28_298 ();
 FILLCELL_X1 FILLER_0_28_302 ();
 FILLCELL_X1 FILLER_0_28_318 ();
 FILLCELL_X2 FILLER_0_28_322 ();
 FILLCELL_X8 FILLER_0_28_327 ();
 FILLCELL_X2 FILLER_0_28_335 ();
 FILLCELL_X4 FILLER_0_28_357 ();
 FILLCELL_X1 FILLER_0_28_361 ();
 FILLCELL_X2 FILLER_0_28_365 ();
 FILLCELL_X1 FILLER_0_28_367 ();
 FILLCELL_X4 FILLER_0_28_372 ();
 FILLCELL_X1 FILLER_0_28_376 ();
 FILLCELL_X4 FILLER_0_28_380 ();
 FILLCELL_X1 FILLER_0_29_1 ();
 FILLCELL_X1 FILLER_0_29_8 ();
 FILLCELL_X1 FILLER_0_29_19 ();
 FILLCELL_X2 FILLER_0_29_52 ();
 FILLCELL_X1 FILLER_0_29_60 ();
 FILLCELL_X1 FILLER_0_29_67 ();
 FILLCELL_X2 FILLER_0_29_71 ();
 FILLCELL_X1 FILLER_0_29_73 ();
 FILLCELL_X1 FILLER_0_29_76 ();
 FILLCELL_X2 FILLER_0_29_80 ();
 FILLCELL_X1 FILLER_0_29_82 ();
 FILLCELL_X2 FILLER_0_29_87 ();
 FILLCELL_X1 FILLER_0_29_89 ();
 FILLCELL_X1 FILLER_0_29_120 ();
 FILLCELL_X1 FILLER_0_29_130 ();
 FILLCELL_X2 FILLER_0_29_134 ();
 FILLCELL_X1 FILLER_0_29_153 ();
 FILLCELL_X4 FILLER_0_29_161 ();
 FILLCELL_X1 FILLER_0_29_165 ();
 FILLCELL_X1 FILLER_0_29_179 ();
 FILLCELL_X1 FILLER_0_29_193 ();
 FILLCELL_X1 FILLER_0_29_203 ();
 FILLCELL_X2 FILLER_0_29_223 ();
 FILLCELL_X1 FILLER_0_29_225 ();
 FILLCELL_X8 FILLER_0_29_236 ();
 FILLCELL_X1 FILLER_0_29_244 ();
 FILLCELL_X2 FILLER_0_29_258 ();
 FILLCELL_X1 FILLER_0_29_266 ();
 FILLCELL_X1 FILLER_0_29_293 ();
 FILLCELL_X2 FILLER_0_29_307 ();
 FILLCELL_X2 FILLER_0_29_315 ();
 FILLCELL_X1 FILLER_0_29_324 ();
 FILLCELL_X1 FILLER_0_29_327 ();
 FILLCELL_X1 FILLER_0_29_331 ();
 FILLCELL_X2 FILLER_0_29_342 ();
 FILLCELL_X1 FILLER_0_29_344 ();
 FILLCELL_X4 FILLER_0_29_351 ();
 FILLCELL_X1 FILLER_0_29_355 ();
 FILLCELL_X8 FILLER_0_29_360 ();
 FILLCELL_X4 FILLER_0_29_368 ();
 FILLCELL_X2 FILLER_0_29_372 ();
 FILLCELL_X1 FILLER_0_29_374 ();
 FILLCELL_X4 FILLER_0_29_382 ();
 FILLCELL_X2 FILLER_0_29_386 ();
 FILLCELL_X4 FILLER_0_30_1 ();
 FILLCELL_X1 FILLER_0_30_5 ();
 FILLCELL_X1 FILLER_0_30_30 ();
 FILLCELL_X1 FILLER_0_30_43 ();
 FILLCELL_X2 FILLER_0_30_50 ();
 FILLCELL_X1 FILLER_0_30_57 ();
 FILLCELL_X2 FILLER_0_30_64 ();
 FILLCELL_X2 FILLER_0_30_70 ();
 FILLCELL_X2 FILLER_0_30_78 ();
 FILLCELL_X1 FILLER_0_30_80 ();
 FILLCELL_X2 FILLER_0_30_87 ();
 FILLCELL_X4 FILLER_0_30_117 ();
 FILLCELL_X2 FILLER_0_30_121 ();
 FILLCELL_X4 FILLER_0_30_133 ();
 FILLCELL_X2 FILLER_0_30_137 ();
 FILLCELL_X1 FILLER_0_30_167 ();
 FILLCELL_X4 FILLER_0_30_174 ();
 FILLCELL_X1 FILLER_0_30_178 ();
 FILLCELL_X4 FILLER_0_30_185 ();
 FILLCELL_X4 FILLER_0_30_203 ();
 FILLCELL_X1 FILLER_0_30_207 ();
 FILLCELL_X4 FILLER_0_30_221 ();
 FILLCELL_X1 FILLER_0_30_225 ();
 FILLCELL_X4 FILLER_0_30_236 ();
 FILLCELL_X2 FILLER_0_30_240 ();
 FILLCELL_X1 FILLER_0_30_242 ();
 FILLCELL_X2 FILLER_0_30_265 ();
 FILLCELL_X1 FILLER_0_30_268 ();
 FILLCELL_X4 FILLER_0_30_282 ();
 FILLCELL_X2 FILLER_0_30_290 ();
 FILLCELL_X1 FILLER_0_30_292 ();
 FILLCELL_X4 FILLER_0_30_365 ();
 FILLCELL_X2 FILLER_0_30_369 ();
 FILLCELL_X2 FILLER_0_31_24 ();
 FILLCELL_X1 FILLER_0_31_26 ();
 FILLCELL_X1 FILLER_0_31_32 ();
 FILLCELL_X8 FILLER_0_31_40 ();
 FILLCELL_X4 FILLER_0_31_48 ();
 FILLCELL_X1 FILLER_0_31_52 ();
 FILLCELL_X4 FILLER_0_31_67 ();
 FILLCELL_X2 FILLER_0_31_71 ();
 FILLCELL_X2 FILLER_0_31_108 ();
 FILLCELL_X8 FILLER_0_31_113 ();
 FILLCELL_X2 FILLER_0_31_121 ();
 FILLCELL_X1 FILLER_0_31_123 ();
 FILLCELL_X2 FILLER_0_31_143 ();
 FILLCELL_X1 FILLER_0_31_145 ();
 FILLCELL_X2 FILLER_0_31_163 ();
 FILLCELL_X8 FILLER_0_31_197 ();
 FILLCELL_X4 FILLER_0_31_205 ();
 FILLCELL_X1 FILLER_0_31_209 ();
 FILLCELL_X4 FILLER_0_31_220 ();
 FILLCELL_X2 FILLER_0_31_224 ();
 FILLCELL_X1 FILLER_0_31_226 ();
 FILLCELL_X1 FILLER_0_31_255 ();
 FILLCELL_X2 FILLER_0_31_262 ();
 FILLCELL_X8 FILLER_0_31_273 ();
 FILLCELL_X1 FILLER_0_31_281 ();
 FILLCELL_X4 FILLER_0_31_286 ();
 FILLCELL_X2 FILLER_0_31_290 ();
 FILLCELL_X2 FILLER_0_31_312 ();
 FILLCELL_X1 FILLER_0_31_328 ();
 FILLCELL_X1 FILLER_0_31_335 ();
 FILLCELL_X1 FILLER_0_31_348 ();
 FILLCELL_X1 FILLER_0_31_355 ();
 FILLCELL_X8 FILLER_0_31_378 ();
 FILLCELL_X2 FILLER_0_31_386 ();
 FILLCELL_X4 FILLER_0_32_1 ();
 FILLCELL_X2 FILLER_0_32_5 ();
 FILLCELL_X4 FILLER_0_32_16 ();
 FILLCELL_X2 FILLER_0_32_20 ();
 FILLCELL_X1 FILLER_0_32_22 ();
 FILLCELL_X1 FILLER_0_32_77 ();
 FILLCELL_X2 FILLER_0_32_96 ();
 FILLCELL_X1 FILLER_0_32_98 ();
 FILLCELL_X8 FILLER_0_32_118 ();
 FILLCELL_X4 FILLER_0_32_126 ();
 FILLCELL_X2 FILLER_0_32_134 ();
 FILLCELL_X1 FILLER_0_32_149 ();
 FILLCELL_X1 FILLER_0_32_153 ();
 FILLCELL_X1 FILLER_0_32_157 ();
 FILLCELL_X1 FILLER_0_32_161 ();
 FILLCELL_X1 FILLER_0_32_168 ();
 FILLCELL_X1 FILLER_0_32_175 ();
 FILLCELL_X2 FILLER_0_32_196 ();
 FILLCELL_X8 FILLER_0_32_201 ();
 FILLCELL_X2 FILLER_0_32_209 ();
 FILLCELL_X1 FILLER_0_32_211 ();
 FILLCELL_X2 FILLER_0_32_221 ();
 FILLCELL_X1 FILLER_0_32_238 ();
 FILLCELL_X2 FILLER_0_32_244 ();
 FILLCELL_X1 FILLER_0_32_251 ();
 FILLCELL_X2 FILLER_0_32_256 ();
 FILLCELL_X4 FILLER_0_32_263 ();
 FILLCELL_X4 FILLER_0_32_268 ();
 FILLCELL_X1 FILLER_0_32_272 ();
 FILLCELL_X1 FILLER_0_32_292 ();
 FILLCELL_X2 FILLER_0_32_320 ();
 FILLCELL_X2 FILLER_0_32_325 ();
 FILLCELL_X1 FILLER_0_32_327 ();
 FILLCELL_X1 FILLER_0_32_334 ();
 FILLCELL_X16 FILLER_0_32_360 ();
 FILLCELL_X8 FILLER_0_32_376 ();
 FILLCELL_X4 FILLER_0_32_384 ();
 FILLCELL_X8 FILLER_0_33_1 ();
 FILLCELL_X2 FILLER_0_33_15 ();
 FILLCELL_X4 FILLER_0_33_21 ();
 FILLCELL_X1 FILLER_0_33_31 ();
 FILLCELL_X2 FILLER_0_33_35 ();
 FILLCELL_X2 FILLER_0_33_39 ();
 FILLCELL_X1 FILLER_0_33_52 ();
 FILLCELL_X4 FILLER_0_33_57 ();
 FILLCELL_X2 FILLER_0_33_61 ();
 FILLCELL_X8 FILLER_0_33_66 ();
 FILLCELL_X2 FILLER_0_33_74 ();
 FILLCELL_X1 FILLER_0_33_76 ();
 FILLCELL_X1 FILLER_0_33_83 ();
 FILLCELL_X4 FILLER_0_33_90 ();
 FILLCELL_X1 FILLER_0_33_114 ();
 FILLCELL_X4 FILLER_0_33_118 ();
 FILLCELL_X2 FILLER_0_33_122 ();
 FILLCELL_X1 FILLER_0_33_124 ();
 FILLCELL_X2 FILLER_0_33_159 ();
 FILLCELL_X2 FILLER_0_33_167 ();
 FILLCELL_X1 FILLER_0_33_169 ();
 FILLCELL_X2 FILLER_0_33_173 ();
 FILLCELL_X4 FILLER_0_33_179 ();
 FILLCELL_X1 FILLER_0_33_183 ();
 FILLCELL_X2 FILLER_0_33_206 ();
 FILLCELL_X1 FILLER_0_33_212 ();
 FILLCELL_X2 FILLER_0_33_217 ();
 FILLCELL_X8 FILLER_0_33_245 ();
 FILLCELL_X1 FILLER_0_33_259 ();
 FILLCELL_X16 FILLER_0_33_266 ();
 FILLCELL_X2 FILLER_0_33_291 ();
 FILLCELL_X4 FILLER_0_33_304 ();
 FILLCELL_X1 FILLER_0_33_308 ();
 FILLCELL_X1 FILLER_0_33_316 ();
 FILLCELL_X2 FILLER_0_33_327 ();
 FILLCELL_X1 FILLER_0_33_343 ();
 FILLCELL_X1 FILLER_0_33_355 ();
 FILLCELL_X16 FILLER_0_33_363 ();
 FILLCELL_X2 FILLER_0_33_379 ();
 FILLCELL_X2 FILLER_0_33_385 ();
 FILLCELL_X1 FILLER_0_33_387 ();
 FILLCELL_X8 FILLER_0_34_1 ();
 FILLCELL_X1 FILLER_0_34_26 ();
 FILLCELL_X1 FILLER_0_34_44 ();
 FILLCELL_X1 FILLER_0_34_55 ();
 FILLCELL_X1 FILLER_0_34_60 ();
 FILLCELL_X2 FILLER_0_34_67 ();
 FILLCELL_X2 FILLER_0_34_72 ();
 FILLCELL_X2 FILLER_0_34_80 ();
 FILLCELL_X1 FILLER_0_34_82 ();
 FILLCELL_X2 FILLER_0_34_86 ();
 FILLCELL_X1 FILLER_0_34_88 ();
 FILLCELL_X4 FILLER_0_34_90 ();
 FILLCELL_X1 FILLER_0_34_94 ();
 FILLCELL_X4 FILLER_0_34_101 ();
 FILLCELL_X2 FILLER_0_34_105 ();
 FILLCELL_X1 FILLER_0_34_107 ();
 FILLCELL_X1 FILLER_0_34_167 ();
 FILLCELL_X1 FILLER_0_34_174 ();
 FILLCELL_X1 FILLER_0_34_185 ();
 FILLCELL_X1 FILLER_0_34_193 ();
 FILLCELL_X1 FILLER_0_34_207 ();
 FILLCELL_X8 FILLER_0_34_214 ();
 FILLCELL_X1 FILLER_0_34_268 ();
 FILLCELL_X1 FILLER_0_34_298 ();
 FILLCELL_X4 FILLER_0_34_325 ();
 FILLCELL_X1 FILLER_0_34_329 ();
 FILLCELL_X2 FILLER_0_34_344 ();
 FILLCELL_X16 FILLER_0_34_361 ();
 FILLCELL_X8 FILLER_0_34_377 ();
 FILLCELL_X2 FILLER_0_34_385 ();
 FILLCELL_X1 FILLER_0_34_387 ();
 FILLCELL_X4 FILLER_0_35_1 ();
 FILLCELL_X1 FILLER_0_35_5 ();
 FILLCELL_X1 FILLER_0_35_26 ();
 FILLCELL_X8 FILLER_0_35_40 ();
 FILLCELL_X2 FILLER_0_35_48 ();
 FILLCELL_X1 FILLER_0_35_50 ();
 FILLCELL_X1 FILLER_0_35_60 ();
 FILLCELL_X4 FILLER_0_35_100 ();
 FILLCELL_X2 FILLER_0_35_104 ();
 FILLCELL_X1 FILLER_0_35_108 ();
 FILLCELL_X8 FILLER_0_35_115 ();
 FILLCELL_X4 FILLER_0_35_154 ();
 FILLCELL_X1 FILLER_0_35_158 ();
 FILLCELL_X1 FILLER_0_35_165 ();
 FILLCELL_X8 FILLER_0_35_168 ();
 FILLCELL_X2 FILLER_0_35_176 ();
 FILLCELL_X4 FILLER_0_35_179 ();
 FILLCELL_X2 FILLER_0_35_183 ();
 FILLCELL_X1 FILLER_0_35_185 ();
 FILLCELL_X1 FILLER_0_35_206 ();
 FILLCELL_X2 FILLER_0_35_211 ();
 FILLCELL_X2 FILLER_0_35_233 ();
 FILLCELL_X2 FILLER_0_35_273 ();
 FILLCELL_X2 FILLER_0_35_292 ();
 FILLCELL_X1 FILLER_0_35_294 ();
 FILLCELL_X2 FILLER_0_35_313 ();
 FILLCELL_X1 FILLER_0_35_315 ();
 FILLCELL_X2 FILLER_0_35_331 ();
 FILLCELL_X1 FILLER_0_35_333 ();
 FILLCELL_X2 FILLER_0_35_340 ();
 FILLCELL_X2 FILLER_0_35_345 ();
 FILLCELL_X2 FILLER_0_35_354 ();
 FILLCELL_X16 FILLER_0_35_363 ();
 FILLCELL_X8 FILLER_0_35_379 ();
 FILLCELL_X1 FILLER_0_35_387 ();
 FILLCELL_X2 FILLER_0_36_1 ();
 FILLCELL_X2 FILLER_0_36_17 ();
 FILLCELL_X1 FILLER_0_36_51 ();
 FILLCELL_X2 FILLER_0_36_75 ();
 FILLCELL_X4 FILLER_0_36_83 ();
 FILLCELL_X2 FILLER_0_36_87 ();
 FILLCELL_X1 FILLER_0_36_97 ();
 FILLCELL_X1 FILLER_0_36_103 ();
 FILLCELL_X1 FILLER_0_36_110 ();
 FILLCELL_X2 FILLER_0_36_116 ();
 FILLCELL_X1 FILLER_0_36_124 ();
 FILLCELL_X2 FILLER_0_36_132 ();
 FILLCELL_X1 FILLER_0_36_153 ();
 FILLCELL_X1 FILLER_0_36_160 ();
 FILLCELL_X1 FILLER_0_36_170 ();
 FILLCELL_X2 FILLER_0_36_175 ();
 FILLCELL_X4 FILLER_0_36_184 ();
 FILLCELL_X4 FILLER_0_36_192 ();
 FILLCELL_X8 FILLER_0_36_215 ();
 FILLCELL_X1 FILLER_0_36_223 ();
 FILLCELL_X2 FILLER_0_36_250 ();
 FILLCELL_X1 FILLER_0_36_261 ();
 FILLCELL_X2 FILLER_0_36_265 ();
 FILLCELL_X4 FILLER_0_36_273 ();
 FILLCELL_X1 FILLER_0_36_277 ();
 FILLCELL_X1 FILLER_0_36_284 ();
 FILLCELL_X2 FILLER_0_36_289 ();
 FILLCELL_X2 FILLER_0_36_324 ();
 FILLCELL_X4 FILLER_0_36_330 ();
 FILLCELL_X4 FILLER_0_36_337 ();
 FILLCELL_X2 FILLER_0_36_347 ();
 FILLCELL_X1 FILLER_0_36_349 ();
 FILLCELL_X1 FILLER_0_36_354 ();
 FILLCELL_X4 FILLER_0_36_361 ();
 FILLCELL_X2 FILLER_0_36_365 ();
 FILLCELL_X1 FILLER_0_36_367 ();
 FILLCELL_X2 FILLER_0_36_385 ();
 FILLCELL_X1 FILLER_0_36_387 ();
 FILLCELL_X4 FILLER_0_37_1 ();
 FILLCELL_X2 FILLER_0_37_5 ();
 FILLCELL_X1 FILLER_0_37_35 ();
 FILLCELL_X1 FILLER_0_37_41 ();
 FILLCELL_X1 FILLER_0_37_45 ();
 FILLCELL_X1 FILLER_0_37_49 ();
 FILLCELL_X2 FILLER_0_37_53 ();
 FILLCELL_X2 FILLER_0_37_58 ();
 FILLCELL_X1 FILLER_0_37_66 ();
 FILLCELL_X2 FILLER_0_37_84 ();
 FILLCELL_X1 FILLER_0_37_86 ();
 FILLCELL_X1 FILLER_0_37_102 ();
 FILLCELL_X1 FILLER_0_37_112 ();
 FILLCELL_X1 FILLER_0_37_149 ();
 FILLCELL_X4 FILLER_0_37_157 ();
 FILLCELL_X1 FILLER_0_37_171 ();
 FILLCELL_X2 FILLER_0_37_176 ();
 FILLCELL_X4 FILLER_0_37_185 ();
 FILLCELL_X1 FILLER_0_37_189 ();
 FILLCELL_X1 FILLER_0_37_193 ();
 FILLCELL_X8 FILLER_0_37_203 ();
 FILLCELL_X2 FILLER_0_37_211 ();
 FILLCELL_X4 FILLER_0_37_255 ();
 FILLCELL_X8 FILLER_0_37_269 ();
 FILLCELL_X2 FILLER_0_37_277 ();
 FILLCELL_X1 FILLER_0_37_279 ();
 FILLCELL_X8 FILLER_0_37_289 ();
 FILLCELL_X2 FILLER_0_37_316 ();
 FILLCELL_X8 FILLER_0_37_340 ();
 FILLCELL_X1 FILLER_0_37_348 ();
 FILLCELL_X1 FILLER_0_37_355 ();
 FILLCELL_X8 FILLER_0_37_357 ();
 FILLCELL_X2 FILLER_0_37_365 ();
 FILLCELL_X1 FILLER_0_37_367 ();
 FILLCELL_X2 FILLER_0_37_385 ();
 FILLCELL_X1 FILLER_0_37_387 ();
 FILLCELL_X4 FILLER_0_38_1 ();
 FILLCELL_X2 FILLER_0_38_11 ();
 FILLCELL_X2 FILLER_0_38_29 ();
 FILLCELL_X1 FILLER_0_38_31 ();
 FILLCELL_X1 FILLER_0_38_55 ();
 FILLCELL_X8 FILLER_0_38_62 ();
 FILLCELL_X2 FILLER_0_38_70 ();
 FILLCELL_X1 FILLER_0_38_72 ();
 FILLCELL_X1 FILLER_0_38_82 ();
 FILLCELL_X4 FILLER_0_38_90 ();
 FILLCELL_X2 FILLER_0_38_94 ();
 FILLCELL_X4 FILLER_0_38_133 ();
 FILLCELL_X1 FILLER_0_38_137 ();
 FILLCELL_X4 FILLER_0_38_140 ();
 FILLCELL_X2 FILLER_0_38_169 ();
 FILLCELL_X1 FILLER_0_38_171 ();
 FILLCELL_X2 FILLER_0_38_178 ();
 FILLCELL_X4 FILLER_0_38_183 ();
 FILLCELL_X2 FILLER_0_38_193 ();
 FILLCELL_X4 FILLER_0_38_201 ();
 FILLCELL_X4 FILLER_0_38_223 ();
 FILLCELL_X1 FILLER_0_38_227 ();
 FILLCELL_X2 FILLER_0_38_254 ();
 FILLCELL_X4 FILLER_0_38_261 ();
 FILLCELL_X2 FILLER_0_38_265 ();
 FILLCELL_X4 FILLER_0_38_278 ();
 FILLCELL_X1 FILLER_0_38_282 ();
 FILLCELL_X1 FILLER_0_38_289 ();
 FILLCELL_X2 FILLER_0_38_293 ();
 FILLCELL_X2 FILLER_0_38_301 ();
 FILLCELL_X2 FILLER_0_38_306 ();
 FILLCELL_X1 FILLER_0_38_308 ();
 FILLCELL_X2 FILLER_0_38_329 ();
 FILLCELL_X8 FILLER_0_38_333 ();
 FILLCELL_X4 FILLER_0_38_341 ();
 FILLCELL_X2 FILLER_0_38_345 ();
 FILLCELL_X32 FILLER_0_38_356 ();
 FILLCELL_X4 FILLER_0_39_1 ();
 FILLCELL_X2 FILLER_0_39_5 ();
 FILLCELL_X4 FILLER_0_39_16 ();
 FILLCELL_X2 FILLER_0_39_45 ();
 FILLCELL_X8 FILLER_0_39_64 ();
 FILLCELL_X2 FILLER_0_39_72 ();
 FILLCELL_X2 FILLER_0_39_91 ();
 FILLCELL_X4 FILLER_0_39_97 ();
 FILLCELL_X4 FILLER_0_39_104 ();
 FILLCELL_X2 FILLER_0_39_108 ();
 FILLCELL_X1 FILLER_0_39_110 ();
 FILLCELL_X2 FILLER_0_39_117 ();
 FILLCELL_X4 FILLER_0_39_125 ();
 FILLCELL_X1 FILLER_0_39_129 ();
 FILLCELL_X4 FILLER_0_39_139 ();
 FILLCELL_X2 FILLER_0_39_143 ();
 FILLCELL_X1 FILLER_0_39_145 ();
 FILLCELL_X1 FILLER_0_39_158 ();
 FILLCELL_X8 FILLER_0_39_162 ();
 FILLCELL_X2 FILLER_0_39_170 ();
 FILLCELL_X2 FILLER_0_39_179 ();
 FILLCELL_X2 FILLER_0_39_187 ();
 FILLCELL_X1 FILLER_0_39_189 ();
 FILLCELL_X2 FILLER_0_39_206 ();
 FILLCELL_X1 FILLER_0_39_208 ();
 FILLCELL_X4 FILLER_0_39_218 ();
 FILLCELL_X1 FILLER_0_39_222 ();
 FILLCELL_X2 FILLER_0_39_227 ();
 FILLCELL_X4 FILLER_0_39_237 ();
 FILLCELL_X1 FILLER_0_39_261 ();
 FILLCELL_X1 FILLER_0_39_297 ();
 FILLCELL_X2 FILLER_0_39_335 ();
 FILLCELL_X1 FILLER_0_39_355 ();
 FILLCELL_X8 FILLER_0_39_363 ();
 FILLCELL_X4 FILLER_0_39_371 ();
 FILLCELL_X1 FILLER_0_39_375 ();
 FILLCELL_X8 FILLER_0_39_380 ();
 FILLCELL_X8 FILLER_0_40_1 ();
 FILLCELL_X2 FILLER_0_40_9 ();
 FILLCELL_X8 FILLER_0_40_14 ();
 FILLCELL_X4 FILLER_0_40_22 ();
 FILLCELL_X1 FILLER_0_40_29 ();
 FILLCELL_X8 FILLER_0_40_39 ();
 FILLCELL_X2 FILLER_0_40_53 ();
 FILLCELL_X4 FILLER_0_40_61 ();
 FILLCELL_X1 FILLER_0_40_90 ();
 FILLCELL_X2 FILLER_0_40_107 ();
 FILLCELL_X1 FILLER_0_40_109 ();
 FILLCELL_X2 FILLER_0_40_116 ();
 FILLCELL_X8 FILLER_0_40_120 ();
 FILLCELL_X2 FILLER_0_40_128 ();
 FILLCELL_X1 FILLER_0_40_130 ();
 FILLCELL_X2 FILLER_0_40_141 ();
 FILLCELL_X1 FILLER_0_40_143 ();
 FILLCELL_X1 FILLER_0_40_150 ();
 FILLCELL_X4 FILLER_0_40_157 ();
 FILLCELL_X1 FILLER_0_40_175 ();
 FILLCELL_X1 FILLER_0_40_179 ();
 FILLCELL_X1 FILLER_0_40_186 ();
 FILLCELL_X1 FILLER_0_40_191 ();
 FILLCELL_X4 FILLER_0_40_207 ();
 FILLCELL_X1 FILLER_0_40_221 ();
 FILLCELL_X1 FILLER_0_40_262 ();
 FILLCELL_X1 FILLER_0_40_268 ();
 FILLCELL_X1 FILLER_0_40_280 ();
 FILLCELL_X1 FILLER_0_40_289 ();
 FILLCELL_X2 FILLER_0_40_301 ();
 FILLCELL_X2 FILLER_0_40_314 ();
 FILLCELL_X1 FILLER_0_40_316 ();
 FILLCELL_X1 FILLER_0_40_320 ();
 FILLCELL_X2 FILLER_0_40_323 ();
 FILLCELL_X4 FILLER_0_40_329 ();
 FILLCELL_X1 FILLER_0_40_333 ();
 FILLCELL_X2 FILLER_0_40_350 ();
 FILLCELL_X1 FILLER_0_40_358 ();
 FILLCELL_X16 FILLER_0_40_365 ();
 FILLCELL_X4 FILLER_0_40_381 ();
 FILLCELL_X2 FILLER_0_40_385 ();
 FILLCELL_X1 FILLER_0_40_387 ();
 FILLCELL_X4 FILLER_0_41_1 ();
 FILLCELL_X2 FILLER_0_41_5 ();
 FILLCELL_X1 FILLER_0_41_7 ();
 FILLCELL_X1 FILLER_0_41_28 ();
 FILLCELL_X1 FILLER_0_41_35 ();
 FILLCELL_X1 FILLER_0_41_40 ();
 FILLCELL_X2 FILLER_0_41_46 ();
 FILLCELL_X1 FILLER_0_41_61 ();
 FILLCELL_X2 FILLER_0_41_77 ();
 FILLCELL_X2 FILLER_0_41_88 ();
 FILLCELL_X4 FILLER_0_41_100 ();
 FILLCELL_X4 FILLER_0_41_127 ();
 FILLCELL_X1 FILLER_0_41_131 ();
 FILLCELL_X2 FILLER_0_41_145 ();
 FILLCELL_X2 FILLER_0_41_150 ();
 FILLCELL_X4 FILLER_0_41_161 ();
 FILLCELL_X2 FILLER_0_41_165 ();
 FILLCELL_X1 FILLER_0_41_167 ();
 FILLCELL_X1 FILLER_0_41_181 ();
 FILLCELL_X4 FILLER_0_41_191 ();
 FILLCELL_X1 FILLER_0_41_195 ();
 FILLCELL_X4 FILLER_0_41_208 ();
 FILLCELL_X8 FILLER_0_41_225 ();
 FILLCELL_X4 FILLER_0_41_233 ();
 FILLCELL_X2 FILLER_0_41_237 ();
 FILLCELL_X8 FILLER_0_41_241 ();
 FILLCELL_X4 FILLER_0_41_249 ();
 FILLCELL_X1 FILLER_0_41_289 ();
 FILLCELL_X1 FILLER_0_41_296 ();
 FILLCELL_X2 FILLER_0_41_301 ();
 FILLCELL_X1 FILLER_0_41_319 ();
 FILLCELL_X1 FILLER_0_41_326 ();
 FILLCELL_X1 FILLER_0_41_339 ();
 FILLCELL_X4 FILLER_0_41_352 ();
 FILLCELL_X16 FILLER_0_41_357 ();
 FILLCELL_X8 FILLER_0_41_373 ();
 FILLCELL_X4 FILLER_0_41_381 ();
 FILLCELL_X2 FILLER_0_41_385 ();
 FILLCELL_X1 FILLER_0_41_387 ();
 FILLCELL_X8 FILLER_0_42_1 ();
 FILLCELL_X2 FILLER_0_42_9 ();
 FILLCELL_X1 FILLER_0_42_11 ();
 FILLCELL_X4 FILLER_0_42_14 ();
 FILLCELL_X2 FILLER_0_42_38 ();
 FILLCELL_X4 FILLER_0_42_54 ();
 FILLCELL_X2 FILLER_0_42_58 ();
 FILLCELL_X1 FILLER_0_42_66 ();
 FILLCELL_X2 FILLER_0_42_80 ();
 FILLCELL_X1 FILLER_0_42_82 ();
 FILLCELL_X2 FILLER_0_42_87 ();
 FILLCELL_X2 FILLER_0_42_99 ();
 FILLCELL_X1 FILLER_0_42_101 ();
 FILLCELL_X4 FILLER_0_42_106 ();
 FILLCELL_X2 FILLER_0_42_110 ();
 FILLCELL_X1 FILLER_0_42_112 ();
 FILLCELL_X1 FILLER_0_42_132 ();
 FILLCELL_X1 FILLER_0_42_142 ();
 FILLCELL_X2 FILLER_0_42_149 ();
 FILLCELL_X1 FILLER_0_42_157 ();
 FILLCELL_X2 FILLER_0_42_162 ();
 FILLCELL_X4 FILLER_0_42_176 ();
 FILLCELL_X2 FILLER_0_42_180 ();
 FILLCELL_X1 FILLER_0_42_182 ();
 FILLCELL_X4 FILLER_0_42_192 ();
 FILLCELL_X4 FILLER_0_42_207 ();
 FILLCELL_X1 FILLER_0_42_211 ();
 FILLCELL_X8 FILLER_0_42_229 ();
 FILLCELL_X4 FILLER_0_42_249 ();
 FILLCELL_X2 FILLER_0_42_253 ();
 FILLCELL_X1 FILLER_0_42_255 ();
 FILLCELL_X2 FILLER_0_42_265 ();
 FILLCELL_X2 FILLER_0_42_284 ();
 FILLCELL_X1 FILLER_0_42_286 ();
 FILLCELL_X1 FILLER_0_42_290 ();
 FILLCELL_X2 FILLER_0_42_297 ();
 FILLCELL_X1 FILLER_0_42_317 ();
 FILLCELL_X2 FILLER_0_42_324 ();
 FILLCELL_X2 FILLER_0_42_329 ();
 FILLCELL_X2 FILLER_0_42_333 ();
 FILLCELL_X1 FILLER_0_42_356 ();
 FILLCELL_X8 FILLER_0_42_363 ();
 FILLCELL_X8 FILLER_0_42_379 ();
 FILLCELL_X1 FILLER_0_42_387 ();
 FILLCELL_X16 FILLER_0_43_1 ();
 FILLCELL_X8 FILLER_0_43_17 ();
 FILLCELL_X4 FILLER_0_43_25 ();
 FILLCELL_X2 FILLER_0_43_29 ();
 FILLCELL_X1 FILLER_0_43_49 ();
 FILLCELL_X2 FILLER_0_43_54 ();
 FILLCELL_X2 FILLER_0_43_62 ();
 FILLCELL_X2 FILLER_0_43_70 ();
 FILLCELL_X2 FILLER_0_43_75 ();
 FILLCELL_X1 FILLER_0_43_77 ();
 FILLCELL_X1 FILLER_0_43_112 ();
 FILLCELL_X8 FILLER_0_43_119 ();
 FILLCELL_X1 FILLER_0_43_127 ();
 FILLCELL_X2 FILLER_0_43_131 ();
 FILLCELL_X2 FILLER_0_43_139 ();
 FILLCELL_X8 FILLER_0_43_145 ();
 FILLCELL_X2 FILLER_0_43_153 ();
 FILLCELL_X2 FILLER_0_43_185 ();
 FILLCELL_X1 FILLER_0_43_206 ();
 FILLCELL_X4 FILLER_0_43_216 ();
 FILLCELL_X4 FILLER_0_43_222 ();
 FILLCELL_X4 FILLER_0_43_228 ();
 FILLCELL_X1 FILLER_0_43_254 ();
 FILLCELL_X2 FILLER_0_43_271 ();
 FILLCELL_X8 FILLER_0_43_277 ();
 FILLCELL_X2 FILLER_0_43_288 ();
 FILLCELL_X4 FILLER_0_43_299 ();
 FILLCELL_X1 FILLER_0_43_306 ();
 FILLCELL_X1 FILLER_0_43_311 ();
 FILLCELL_X2 FILLER_0_43_322 ();
 FILLCELL_X1 FILLER_0_43_324 ();
 FILLCELL_X1 FILLER_0_43_357 ();
 FILLCELL_X1 FILLER_0_43_362 ();
 FILLCELL_X1 FILLER_0_43_369 ();
 FILLCELL_X1 FILLER_0_43_374 ();
 FILLCELL_X8 FILLER_0_43_380 ();
 FILLCELL_X16 FILLER_0_44_1 ();
 FILLCELL_X8 FILLER_0_44_17 ();
 FILLCELL_X2 FILLER_0_44_40 ();
 FILLCELL_X8 FILLER_0_44_48 ();
 FILLCELL_X2 FILLER_0_44_56 ();
 FILLCELL_X8 FILLER_0_44_73 ();
 FILLCELL_X2 FILLER_0_44_81 ();
 FILLCELL_X1 FILLER_0_44_94 ();
 FILLCELL_X2 FILLER_0_44_101 ();
 FILLCELL_X2 FILLER_0_44_105 ();
 FILLCELL_X2 FILLER_0_44_110 ();
 FILLCELL_X8 FILLER_0_44_121 ();
 FILLCELL_X2 FILLER_0_44_129 ();
 FILLCELL_X16 FILLER_0_44_140 ();
 FILLCELL_X1 FILLER_0_44_156 ();
 FILLCELL_X1 FILLER_0_44_166 ();
 FILLCELL_X1 FILLER_0_44_171 ();
 FILLCELL_X1 FILLER_0_44_176 ();
 FILLCELL_X1 FILLER_0_44_183 ();
 FILLCELL_X1 FILLER_0_44_189 ();
 FILLCELL_X1 FILLER_0_44_193 ();
 FILLCELL_X1 FILLER_0_44_201 ();
 FILLCELL_X2 FILLER_0_44_208 ();
 FILLCELL_X1 FILLER_0_44_210 ();
 FILLCELL_X1 FILLER_0_44_215 ();
 FILLCELL_X2 FILLER_0_44_224 ();
 FILLCELL_X1 FILLER_0_44_231 ();
 FILLCELL_X1 FILLER_0_44_261 ();
 FILLCELL_X1 FILLER_0_44_266 ();
 FILLCELL_X1 FILLER_0_44_277 ();
 FILLCELL_X2 FILLER_0_44_315 ();
 FILLCELL_X1 FILLER_0_44_317 ();
 FILLCELL_X1 FILLER_0_44_328 ();
 FILLCELL_X2 FILLER_0_44_331 ();
 FILLCELL_X2 FILLER_0_44_339 ();
 FILLCELL_X2 FILLER_0_44_345 ();
 FILLCELL_X1 FILLER_0_44_347 ();
 FILLCELL_X1 FILLER_0_44_355 ();
 FILLCELL_X1 FILLER_0_44_358 ();
 FILLCELL_X1 FILLER_0_44_371 ();
 FILLCELL_X8 FILLER_0_44_376 ();
 FILLCELL_X4 FILLER_0_44_384 ();
 FILLCELL_X16 FILLER_0_45_1 ();
 FILLCELL_X8 FILLER_0_45_17 ();
 FILLCELL_X1 FILLER_0_45_36 ();
 FILLCELL_X4 FILLER_0_45_41 ();
 FILLCELL_X2 FILLER_0_45_45 ();
 FILLCELL_X1 FILLER_0_45_47 ();
 FILLCELL_X4 FILLER_0_45_65 ();
 FILLCELL_X1 FILLER_0_45_69 ();
 FILLCELL_X2 FILLER_0_45_90 ();
 FILLCELL_X1 FILLER_0_45_95 ();
 FILLCELL_X8 FILLER_0_45_99 ();
 FILLCELL_X4 FILLER_0_45_107 ();
 FILLCELL_X1 FILLER_0_45_111 ();
 FILLCELL_X4 FILLER_0_45_142 ();
 FILLCELL_X2 FILLER_0_45_146 ();
 FILLCELL_X2 FILLER_0_45_154 ();
 FILLCELL_X1 FILLER_0_45_177 ();
 FILLCELL_X2 FILLER_0_45_185 ();
 FILLCELL_X8 FILLER_0_45_205 ();
 FILLCELL_X4 FILLER_0_45_213 ();
 FILLCELL_X1 FILLER_0_45_217 ();
 FILLCELL_X2 FILLER_0_45_224 ();
 FILLCELL_X4 FILLER_0_45_232 ();
 FILLCELL_X1 FILLER_0_45_242 ();
 FILLCELL_X2 FILLER_0_45_245 ();
 FILLCELL_X1 FILLER_0_45_250 ();
 FILLCELL_X2 FILLER_0_45_255 ();
 FILLCELL_X1 FILLER_0_45_261 ();
 FILLCELL_X1 FILLER_0_45_266 ();
 FILLCELL_X1 FILLER_0_45_272 ();
 FILLCELL_X2 FILLER_0_45_279 ();
 FILLCELL_X8 FILLER_0_45_284 ();
 FILLCELL_X1 FILLER_0_45_301 ();
 FILLCELL_X1 FILLER_0_45_305 ();
 FILLCELL_X1 FILLER_0_45_312 ();
 FILLCELL_X2 FILLER_0_45_322 ();
 FILLCELL_X4 FILLER_0_45_333 ();
 FILLCELL_X2 FILLER_0_45_337 ();
 FILLCELL_X1 FILLER_0_45_339 ();
 FILLCELL_X4 FILLER_0_45_346 ();
 FILLCELL_X2 FILLER_0_45_357 ();
 FILLCELL_X16 FILLER_0_46_1 ();
 FILLCELL_X4 FILLER_0_46_17 ();
 FILLCELL_X1 FILLER_0_46_21 ();
 FILLCELL_X4 FILLER_0_46_59 ();
 FILLCELL_X2 FILLER_0_46_63 ();
 FILLCELL_X1 FILLER_0_46_88 ();
 FILLCELL_X4 FILLER_0_46_90 ();
 FILLCELL_X2 FILLER_0_46_94 ();
 FILLCELL_X2 FILLER_0_46_102 ();
 FILLCELL_X2 FILLER_0_46_107 ();
 FILLCELL_X1 FILLER_0_46_128 ();
 FILLCELL_X1 FILLER_0_46_135 ();
 FILLCELL_X1 FILLER_0_46_141 ();
 FILLCELL_X2 FILLER_0_46_144 ();
 FILLCELL_X1 FILLER_0_46_163 ();
 FILLCELL_X2 FILLER_0_46_179 ();
 FILLCELL_X1 FILLER_0_46_181 ();
 FILLCELL_X16 FILLER_0_46_203 ();
 FILLCELL_X8 FILLER_0_46_219 ();
 FILLCELL_X2 FILLER_0_46_250 ();
 FILLCELL_X1 FILLER_0_46_266 ();
 FILLCELL_X2 FILLER_0_46_300 ();
 FILLCELL_X2 FILLER_0_46_311 ();
 FILLCELL_X1 FILLER_0_46_313 ();
 FILLCELL_X2 FILLER_0_46_323 ();
 FILLCELL_X1 FILLER_0_46_331 ();
 FILLCELL_X1 FILLER_0_46_336 ();
 FILLCELL_X2 FILLER_0_46_356 ();
 FILLCELL_X16 FILLER_0_46_367 ();
 FILLCELL_X4 FILLER_0_46_383 ();
 FILLCELL_X1 FILLER_0_46_387 ();
 FILLCELL_X8 FILLER_0_47_1 ();
 FILLCELL_X2 FILLER_0_47_9 ();
 FILLCELL_X1 FILLER_0_47_11 ();
 FILLCELL_X1 FILLER_0_47_32 ();
 FILLCELL_X4 FILLER_0_47_37 ();
 FILLCELL_X2 FILLER_0_47_41 ();
 FILLCELL_X1 FILLER_0_47_48 ();
 FILLCELL_X1 FILLER_0_47_52 ();
 FILLCELL_X1 FILLER_0_47_87 ();
 FILLCELL_X1 FILLER_0_47_124 ();
 FILLCELL_X2 FILLER_0_47_144 ();
 FILLCELL_X1 FILLER_0_47_149 ();
 FILLCELL_X2 FILLER_0_47_176 ();
 FILLCELL_X2 FILLER_0_47_186 ();
 FILLCELL_X1 FILLER_0_47_188 ();
 FILLCELL_X2 FILLER_0_47_203 ();
 FILLCELL_X1 FILLER_0_47_205 ();
 FILLCELL_X1 FILLER_0_47_238 ();
 FILLCELL_X2 FILLER_0_47_249 ();
 FILLCELL_X2 FILLER_0_47_255 ();
 FILLCELL_X2 FILLER_0_47_279 ();
 FILLCELL_X1 FILLER_0_47_281 ();
 FILLCELL_X8 FILLER_0_47_292 ();
 FILLCELL_X4 FILLER_0_47_310 ();
 FILLCELL_X1 FILLER_0_47_349 ();
 FILLCELL_X1 FILLER_0_47_357 ();
 FILLCELL_X1 FILLER_0_47_367 ();
 FILLCELL_X1 FILLER_0_47_372 ();
 FILLCELL_X2 FILLER_0_47_377 ();
 FILLCELL_X4 FILLER_0_47_381 ();
 FILLCELL_X2 FILLER_0_47_385 ();
 FILLCELL_X1 FILLER_0_47_387 ();
 FILLCELL_X16 FILLER_0_48_1 ();
 FILLCELL_X8 FILLER_0_48_17 ();
 FILLCELL_X1 FILLER_0_48_25 ();
 FILLCELL_X1 FILLER_0_48_66 ();
 FILLCELL_X1 FILLER_0_48_83 ();
 FILLCELL_X1 FILLER_0_48_88 ();
 FILLCELL_X1 FILLER_0_48_90 ();
 FILLCELL_X1 FILLER_0_48_103 ();
 FILLCELL_X2 FILLER_0_48_113 ();
 FILLCELL_X2 FILLER_0_48_118 ();
 FILLCELL_X1 FILLER_0_48_136 ();
 FILLCELL_X1 FILLER_0_48_139 ();
 FILLCELL_X1 FILLER_0_48_157 ();
 FILLCELL_X1 FILLER_0_48_162 ();
 FILLCELL_X4 FILLER_0_48_182 ();
 FILLCELL_X4 FILLER_0_48_189 ();
 FILLCELL_X2 FILLER_0_48_193 ();
 FILLCELL_X1 FILLER_0_48_195 ();
 FILLCELL_X4 FILLER_0_48_206 ();
 FILLCELL_X1 FILLER_0_48_210 ();
 FILLCELL_X1 FILLER_0_48_216 ();
 FILLCELL_X2 FILLER_0_48_234 ();
 FILLCELL_X4 FILLER_0_48_263 ();
 FILLCELL_X1 FILLER_0_48_285 ();
 FILLCELL_X1 FILLER_0_48_292 ();
 FILLCELL_X1 FILLER_0_48_302 ();
 FILLCELL_X4 FILLER_0_48_309 ();
 FILLCELL_X2 FILLER_0_48_313 ();
 FILLCELL_X1 FILLER_0_48_315 ();
 FILLCELL_X1 FILLER_0_48_329 ();
 FILLCELL_X4 FILLER_0_48_336 ();
 FILLCELL_X2 FILLER_0_48_354 ();
 FILLCELL_X1 FILLER_0_48_367 ();
 FILLCELL_X2 FILLER_0_48_372 ();
 FILLCELL_X8 FILLER_0_48_380 ();
 FILLCELL_X16 FILLER_0_49_1 ();
 FILLCELL_X8 FILLER_0_49_17 ();
 FILLCELL_X2 FILLER_0_49_25 ();
 FILLCELL_X1 FILLER_0_49_27 ();
 FILLCELL_X2 FILLER_0_49_45 ();
 FILLCELL_X1 FILLER_0_49_63 ();
 FILLCELL_X2 FILLER_0_49_92 ();
 FILLCELL_X2 FILLER_0_49_116 ();
 FILLCELL_X1 FILLER_0_49_128 ();
 FILLCELL_X1 FILLER_0_49_135 ();
 FILLCELL_X1 FILLER_0_49_139 ();
 FILLCELL_X2 FILLER_0_49_146 ();
 FILLCELL_X2 FILLER_0_49_157 ();
 FILLCELL_X1 FILLER_0_49_159 ();
 FILLCELL_X1 FILLER_0_49_199 ();
 FILLCELL_X1 FILLER_0_49_213 ();
 FILLCELL_X1 FILLER_0_49_218 ();
 FILLCELL_X1 FILLER_0_49_223 ();
 FILLCELL_X1 FILLER_0_49_228 ();
 FILLCELL_X1 FILLER_0_49_233 ();
 FILLCELL_X1 FILLER_0_49_243 ();
 FILLCELL_X2 FILLER_0_49_248 ();
 FILLCELL_X4 FILLER_0_49_254 ();
 FILLCELL_X1 FILLER_0_49_270 ();
 FILLCELL_X1 FILLER_0_49_274 ();
 FILLCELL_X1 FILLER_0_49_279 ();
 FILLCELL_X2 FILLER_0_49_286 ();
 FILLCELL_X1 FILLER_0_49_294 ();
 FILLCELL_X2 FILLER_0_49_312 ();
 FILLCELL_X1 FILLER_0_49_323 ();
 FILLCELL_X8 FILLER_0_49_328 ();
 FILLCELL_X2 FILLER_0_49_336 ();
 FILLCELL_X1 FILLER_0_49_355 ();
 FILLCELL_X8 FILLER_0_49_379 ();
 FILLCELL_X1 FILLER_0_49_387 ();
 FILLCELL_X16 FILLER_0_50_1 ();
 FILLCELL_X4 FILLER_0_50_17 ();
 FILLCELL_X1 FILLER_0_50_21 ();
 FILLCELL_X4 FILLER_0_50_43 ();
 FILLCELL_X4 FILLER_0_50_53 ();
 FILLCELL_X2 FILLER_0_50_57 ();
 FILLCELL_X2 FILLER_0_50_73 ();
 FILLCELL_X1 FILLER_0_50_75 ();
 FILLCELL_X2 FILLER_0_50_79 ();
 FILLCELL_X1 FILLER_0_50_81 ();
 FILLCELL_X1 FILLER_0_50_85 ();
 FILLCELL_X1 FILLER_0_50_104 ();
 FILLCELL_X2 FILLER_0_50_111 ();
 FILLCELL_X1 FILLER_0_50_122 ();
 FILLCELL_X2 FILLER_0_50_134 ();
 FILLCELL_X1 FILLER_0_50_136 ();
 FILLCELL_X4 FILLER_0_50_158 ();
 FILLCELL_X1 FILLER_0_50_162 ();
 FILLCELL_X1 FILLER_0_50_172 ();
 FILLCELL_X2 FILLER_0_50_177 ();
 FILLCELL_X1 FILLER_0_50_179 ();
 FILLCELL_X2 FILLER_0_50_184 ();
 FILLCELL_X4 FILLER_0_50_203 ();
 FILLCELL_X1 FILLER_0_50_211 ();
 FILLCELL_X1 FILLER_0_50_223 ();
 FILLCELL_X1 FILLER_0_50_264 ();
 FILLCELL_X1 FILLER_0_50_280 ();
 FILLCELL_X1 FILLER_0_50_285 ();
 FILLCELL_X1 FILLER_0_50_309 ();
 FILLCELL_X1 FILLER_0_50_316 ();
 FILLCELL_X1 FILLER_0_50_321 ();
 FILLCELL_X16 FILLER_0_50_326 ();
 FILLCELL_X4 FILLER_0_50_384 ();
 FILLCELL_X16 FILLER_0_51_1 ();
 FILLCELL_X8 FILLER_0_51_17 ();
 FILLCELL_X4 FILLER_0_51_25 ();
 FILLCELL_X2 FILLER_0_51_29 ();
 FILLCELL_X1 FILLER_0_51_42 ();
 FILLCELL_X1 FILLER_0_51_50 ();
 FILLCELL_X2 FILLER_0_51_54 ();
 FILLCELL_X1 FILLER_0_51_56 ();
 FILLCELL_X1 FILLER_0_51_74 ();
 FILLCELL_X4 FILLER_0_51_81 ();
 FILLCELL_X4 FILLER_0_51_90 ();
 FILLCELL_X2 FILLER_0_51_94 ();
 FILLCELL_X8 FILLER_0_51_101 ();
 FILLCELL_X1 FILLER_0_51_109 ();
 FILLCELL_X2 FILLER_0_51_121 ();
 FILLCELL_X1 FILLER_0_51_126 ();
 FILLCELL_X1 FILLER_0_51_138 ();
 FILLCELL_X2 FILLER_0_51_142 ();
 FILLCELL_X1 FILLER_0_51_144 ();
 FILLCELL_X8 FILLER_0_51_162 ();
 FILLCELL_X2 FILLER_0_51_170 ();
 FILLCELL_X2 FILLER_0_51_179 ();
 FILLCELL_X2 FILLER_0_51_184 ();
 FILLCELL_X1 FILLER_0_51_186 ();
 FILLCELL_X2 FILLER_0_51_198 ();
 FILLCELL_X1 FILLER_0_51_206 ();
 FILLCELL_X1 FILLER_0_51_214 ();
 FILLCELL_X1 FILLER_0_51_218 ();
 FILLCELL_X2 FILLER_0_51_227 ();
 FILLCELL_X16 FILLER_0_51_235 ();
 FILLCELL_X8 FILLER_0_51_251 ();
 FILLCELL_X2 FILLER_0_51_268 ();
 FILLCELL_X2 FILLER_0_51_285 ();
 FILLCELL_X8 FILLER_0_51_298 ();
 FILLCELL_X4 FILLER_0_51_306 ();
 FILLCELL_X1 FILLER_0_51_310 ();
 FILLCELL_X4 FILLER_0_51_314 ();
 FILLCELL_X2 FILLER_0_51_318 ();
 FILLCELL_X1 FILLER_0_51_320 ();
 FILLCELL_X16 FILLER_0_51_338 ();
 FILLCELL_X2 FILLER_0_51_354 ();
 FILLCELL_X4 FILLER_0_51_357 ();
 FILLCELL_X2 FILLER_0_51_361 ();
 FILLCELL_X1 FILLER_0_51_363 ();
 FILLCELL_X1 FILLER_0_51_368 ();
 FILLCELL_X8 FILLER_0_51_376 ();
 FILLCELL_X4 FILLER_0_51_384 ();
endmodule
